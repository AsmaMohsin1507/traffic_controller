// This is the unpowered netlist.
module tiny_user_project (io_in,
    io_oeb,
    io_out);
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire net15;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net16;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net17;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net53;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net54;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net55;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire \mod.cnter_enb_ovf_i1.cnt_val[0] ;
 wire \mod.cnter_enb_ovf_i1.cnt_val[1] ;
 wire \mod.cnter_enb_ovf_i1.cnt_val[2] ;
 wire \mod.cnter_enb_ovf_i1.cnt_val[3] ;
 wire \mod.cnter_enb_ovf_i1.cnt_val[4] ;
 wire \mod.cnter_enb_ovf_i1.overflow ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[0] ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[1] ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[2] ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[3] ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[4] ;
 wire \mod.traffic_sm_inst.traffic_state[0] ;
 wire \mod.traffic_sm_inst.traffic_state[1] ;
 wire \mod.traffic_sm_inst.traffic_state[2] ;
 wire \mod.traffic_sm_inst.traffic_state[3] ;
 wire \mod.traffic_sm_inst.traffic_state[4] ;
 wire \mod.traffic_sm_inst.traffic_state[5] ;
 wire \mod.traffic_sm_inst.traffic_state[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;

 sky130_fd_sc_hd__or3b_1 _067_ (.A(\mod.traffic_sm_inst.traffic_state[5] ),
    .B(\mod.traffic_sm_inst.traffic_state[4] ),
    .C_N(\mod.traffic_sm_inst.traffic_state[6] ),
    .X(_027_));
 sky130_fd_sc_hd__or3b_1 _068_ (.A(\mod.traffic_sm_inst.traffic_state[5] ),
    .B(\mod.traffic_sm_inst.traffic_state[6] ),
    .C_N(\mod.traffic_sm_inst.traffic_state[4] ),
    .X(_028_));
 sky130_fd_sc_hd__nor4_1 _069_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(\mod.traffic_sm_inst.traffic_state[1] ),
    .C(\mod.traffic_sm_inst.traffic_state[3] ),
    .D(\mod.traffic_sm_inst.traffic_state[2] ),
    .Y(_029_));
 sky130_fd_sc_hd__a21boi_4 _070_ (.A1(_027_),
    .A2(_028_),
    .B1_N(_029_),
    .Y(net8));
 sky130_fd_sc_hd__and4bb_1 _071_ (.A_N(\mod.traffic_sm_inst.traffic_state[4] ),
    .B_N(\mod.traffic_sm_inst.traffic_state[6] ),
    .C(_029_),
    .D(\mod.traffic_sm_inst.traffic_state[5] ),
    .X(_030_));
 sky130_fd_sc_hd__clkbuf_2 _072_ (.A(_030_),
    .X(net9));
 sky130_fd_sc_hd__nor2_1 _073_ (.A(net8),
    .B(net9),
    .Y(net7));
 sky130_fd_sc_hd__or4b_1 _074_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(\mod.traffic_sm_inst.traffic_state[1] ),
    .C(\mod.traffic_sm_inst.traffic_state[2] ),
    .D_N(\mod.traffic_sm_inst.traffic_state[3] ),
    .X(_031_));
 sky130_fd_sc_hd__or4b_2 _075_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(\mod.traffic_sm_inst.traffic_state[3] ),
    .C(\mod.traffic_sm_inst.traffic_state[2] ),
    .D_N(\mod.traffic_sm_inst.traffic_state[1] ),
    .X(_032_));
 sky130_fd_sc_hd__or3_1 _076_ (.A(\mod.traffic_sm_inst.traffic_state[5] ),
    .B(\mod.traffic_sm_inst.traffic_state[4] ),
    .C(\mod.traffic_sm_inst.traffic_state[6] ),
    .X(_033_));
 sky130_fd_sc_hd__clkbuf_2 _077_ (.A(_033_),
    .X(_034_));
 sky130_fd_sc_hd__a21oi_2 _078_ (.A1(_031_),
    .A2(_032_),
    .B1(_034_),
    .Y(net5));
 sky130_fd_sc_hd__or4b_1 _079_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(\mod.traffic_sm_inst.traffic_state[1] ),
    .C(\mod.traffic_sm_inst.traffic_state[3] ),
    .D_N(\mod.traffic_sm_inst.traffic_state[2] ),
    .X(_035_));
 sky130_fd_sc_hd__nor2_2 _080_ (.A(_034_),
    .B(_035_),
    .Y(net6));
 sky130_fd_sc_hd__nor2_1 _081_ (.A(net5),
    .B(net6),
    .Y(net4));
 sky130_fd_sc_hd__and4bb_1 _082_ (.A_N(\mod.traffic_sm_inst.traffic_state[5] ),
    .B_N(\mod.traffic_sm_inst.traffic_state[4] ),
    .C(\mod.traffic_sm_inst.traffic_state[6] ),
    .D(_029_),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _083_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .X(_037_));
 sky130_fd_sc_hd__and2b_1 _084_ (.A_N(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .X(_038_));
 sky130_fd_sc_hd__and3_1 _085_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .B(_037_),
    .C(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nor4_1 _086_ (.A(net8),
    .B(net9),
    .C(net5),
    .D(net6),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_1 _087_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(net1),
    .Y(_041_));
 sky130_fd_sc_hd__or3_1 _088_ (.A(\mod.traffic_sm_inst.traffic_state[1] ),
    .B(\mod.traffic_sm_inst.traffic_state[3] ),
    .C(\mod.traffic_sm_inst.traffic_state[2] ),
    .X(_042_));
 sky130_fd_sc_hd__or3_1 _089_ (.A(_034_),
    .B(_041_),
    .C(_042_),
    .X(_043_));
 sky130_fd_sc_hd__a22o_1 _090_ (.A1(_036_),
    .A2(_039_),
    .B1(_040_),
    .B2(_043_),
    .X(_011_));
 sky130_fd_sc_hd__nor2_1 _091_ (.A(_034_),
    .B(_032_),
    .Y(_044_));
 sky130_fd_sc_hd__or3b_1 _092_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .C_N(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .X(_045_));
 sky130_fd_sc_hd__or3_1 _093_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .C(_045_),
    .X(_046_));
 sky130_fd_sc_hd__a21bo_1 _094_ (.A1(_044_),
    .A2(_046_),
    .B1_N(_043_),
    .X(_012_));
 sky130_fd_sc_hd__and2b_1 _095_ (.A_N(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .B(_037_),
    .X(_047_));
 sky130_fd_sc_hd__a21bo_1 _096_ (.A1(_038_),
    .A2(_047_),
    .B1_N(net6),
    .X(_048_));
 sky130_fd_sc_hd__o31ai_1 _097_ (.A1(_034_),
    .A2(_032_),
    .A3(_046_),
    .B1(_048_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _098_ (.A(_045_),
    .Y(_049_));
 sky130_fd_sc_hd__nand3_1 _099_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .C(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__nor2_1 _100_ (.A(_034_),
    .B(_031_),
    .Y(_051_));
 sky130_fd_sc_hd__a32o_1 _101_ (.A1(net6),
    .A2(_038_),
    .A3(_047_),
    .B1(_050_),
    .B2(_051_),
    .X(_014_));
 sky130_fd_sc_hd__and3_1 _102_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .C(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .X(_052_));
 sky130_fd_sc_hd__nand2_1 _103_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .B(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__and4bb_1 _104_ (.A_N(\mod.traffic_sm_inst.traffic_state[5] ),
    .B_N(\mod.traffic_sm_inst.traffic_state[6] ),
    .C(_029_),
    .D(\mod.traffic_sm_inst.traffic_state[4] ),
    .X(_054_));
 sky130_fd_sc_hd__o21a_1 _105_ (.A1(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .A2(_053_),
    .B1(_054_),
    .X(_055_));
 sky130_fd_sc_hd__a41o_1 _106_ (.A1(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .A2(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .A3(_051_),
    .A4(_049_),
    .B1(_055_),
    .X(_015_));
 sky130_fd_sc_hd__nor2_1 _107_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .B(_053_),
    .Y(_056_));
 sky130_fd_sc_hd__and4b_1 _108_ (.A_N(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .C(_038_),
    .D(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .X(_057_));
 sky130_fd_sc_hd__and2b_1 _109_ (.A_N(_057_),
    .B(net9),
    .X(_058_));
 sky130_fd_sc_hd__a21o_1 _110_ (.A1(_054_),
    .A2(_056_),
    .B1(_058_),
    .X(_016_));
 sky130_fd_sc_hd__inv_2 _111_ (.A(_039_),
    .Y(_059_));
 sky130_fd_sc_hd__a22o_1 _112_ (.A1(_036_),
    .A2(_059_),
    .B1(_057_),
    .B2(net9),
    .X(_017_));
 sky130_fd_sc_hd__nor2_1 _113_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[3] ),
    .B(\mod.cnter_enb_ovf_i1.cnt_val[4] ),
    .Y(_060_));
 sky130_fd_sc_hd__and2_1 _114_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i1.cnt_val[0] ),
    .X(_061_));
 sky130_fd_sc_hd__o41a_1 _115_ (.A1(net8),
    .A2(net9),
    .A3(net5),
    .A4(net6),
    .B1(_061_),
    .X(_062_));
 sky130_fd_sc_hd__and3b_1 _116_ (.A_N(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .B(_060_),
    .C(_062_),
    .X(_063_));
 sky130_fd_sc_hd__clkbuf_1 _117_ (.A(_063_),
    .X(_000_));
 sky130_fd_sc_hd__xor2_1 _118_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .B(\mod.cnter_enb_ovf_i1.overflow ),
    .X(_006_));
 sky130_fd_sc_hd__a21oi_1 _119_ (.A1(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .A2(\mod.cnter_enb_ovf_i1.overflow ),
    .B1(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .Y(_064_));
 sky130_fd_sc_hd__and3_1 _120_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .C(\mod.cnter_enb_ovf_i1.overflow ),
    .X(_065_));
 sky130_fd_sc_hd__nor2_1 _121_ (.A(_064_),
    .B(_065_),
    .Y(_007_));
 sky130_fd_sc_hd__and2_1 _122_ (.A(\mod.cnter_enb_ovf_i1.overflow ),
    .B(_052_),
    .X(_066_));
 sky130_fd_sc_hd__nor2_1 _123_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .B(_065_),
    .Y(_018_));
 sky130_fd_sc_hd__a211oi_1 _124_ (.A1(\mod.cnter_enb_ovf_i1.overflow ),
    .A2(_039_),
    .B1(_066_),
    .C1(_018_),
    .Y(_008_));
 sky130_fd_sc_hd__a22oi_1 _125_ (.A1(\mod.cnter_enb_ovf_i1.overflow ),
    .A2(_039_),
    .B1(_066_),
    .B2(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .Y(_019_));
 sky130_fd_sc_hd__o21a_1 _126_ (.A1(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .A2(_066_),
    .B1(_019_),
    .X(_009_));
 sky130_fd_sc_hd__a22o_1 _127_ (.A1(\mod.cnter_enb_ovf_i1.overflow ),
    .A2(_056_),
    .B1(_019_),
    .B2(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .X(_010_));
 sky130_fd_sc_hd__xnor2_1 _128_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[0] ),
    .B(_040_),
    .Y(_001_));
 sky130_fd_sc_hd__o41a_1 _129_ (.A1(net8),
    .A2(net9),
    .A3(net5),
    .A4(net6),
    .B1(\mod.cnter_enb_ovf_i1.cnt_val[0] ),
    .X(_020_));
 sky130_fd_sc_hd__xor2_1 _130_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[1] ),
    .B(_020_),
    .X(_002_));
 sky130_fd_sc_hd__nor2_1 _131_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .B(_060_),
    .Y(_021_));
 sky130_fd_sc_hd__mux2_1 _132_ (.A0(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .A1(_021_),
    .S(_062_),
    .X(_022_));
 sky130_fd_sc_hd__clkbuf_1 _133_ (.A(_022_),
    .X(_003_));
 sky130_fd_sc_hd__xor2_1 _134_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[3] ),
    .B(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _135_ (.A0(\mod.cnter_enb_ovf_i1.cnt_val[3] ),
    .A1(_023_),
    .S(_062_),
    .X(_024_));
 sky130_fd_sc_hd__clkbuf_1 _136_ (.A(_024_),
    .X(_004_));
 sky130_fd_sc_hd__and3_1 _137_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[3] ),
    .B(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .C(_061_),
    .X(_025_));
 sky130_fd_sc_hd__o41a_1 _138_ (.A1(net8),
    .A2(net9),
    .A3(net5),
    .A4(net6),
    .B1(_025_),
    .X(_026_));
 sky130_fd_sc_hd__xor2_1 _139_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[4] ),
    .B(_026_),
    .X(_005_));
 sky130_fd_sc_hd__dfrtp_1 _140_ (.CLK(net12),
    .D(_006_),
    .RESET_B(net10),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[0] ));
 sky130_fd_sc_hd__dfrtp_1 _141_ (.CLK(net13),
    .D(_007_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[1] ));
 sky130_fd_sc_hd__dfrtp_1 _142_ (.CLK(net13),
    .D(_008_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[2] ));
 sky130_fd_sc_hd__dfrtp_1 _143_ (.CLK(net13),
    .D(_009_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[3] ));
 sky130_fd_sc_hd__dfrtp_1 _144_ (.CLK(net12),
    .D(_010_),
    .RESET_B(net10),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[4] ));
 sky130_fd_sc_hd__dfstp_1 _145_ (.CLK(net12),
    .D(_011_),
    .SET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _146_ (.CLK(net12),
    .D(_012_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _147_ (.CLK(net12),
    .D(_013_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _148_ (.CLK(net12),
    .D(_014_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _149_ (.CLK(net12),
    .D(_015_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _150_ (.CLK(net12),
    .D(_016_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _151_ (.CLK(net13),
    .D(_017_),
    .RESET_B(net11),
    .Q(\mod.traffic_sm_inst.traffic_state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _152_ (.CLK(net12),
    .D(_001_),
    .RESET_B(net10),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[0] ));
 sky130_fd_sc_hd__dfrtp_1 _153_ (.CLK(net13),
    .D(_002_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[1] ));
 sky130_fd_sc_hd__dfrtp_1 _154_ (.CLK(net13),
    .D(_003_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[2] ));
 sky130_fd_sc_hd__dfrtp_1 _155_ (.CLK(net13),
    .D(_004_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[3] ));
 sky130_fd_sc_hd__dfrtp_1 _156_ (.CLK(net12),
    .D(_005_),
    .RESET_B(net10),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[4] ));
 sky130_fd_sc_hd__dfrtp_2 _157_ (.CLK(net13),
    .D(_000_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i1.overflow ));
 sky130_fd_sc_hd__conb_1 tiny_user_project_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 tiny_user_project_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 tiny_user_project_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 tiny_user_project_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 tiny_user_project_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 tiny_user_project_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 tiny_user_project_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 tiny_user_project_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 tiny_user_project_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 tiny_user_project_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 tiny_user_project_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 tiny_user_project_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 tiny_user_project_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 tiny_user_project_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 tiny_user_project_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 tiny_user_project_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 tiny_user_project_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 tiny_user_project_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 tiny_user_project_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 tiny_user_project_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 tiny_user_project_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 tiny_user_project_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 tiny_user_project_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 tiny_user_project_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 tiny_user_project_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 tiny_user_project_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 tiny_user_project_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 tiny_user_project_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 tiny_user_project_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 tiny_user_project_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 tiny_user_project_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 tiny_user_project_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 tiny_user_project_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 tiny_user_project_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 tiny_user_project_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 tiny_user_project_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 tiny_user_project_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 tiny_user_project_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 tiny_user_project_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 tiny_user_project_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 tiny_user_project_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 tiny_user_project_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 tiny_user_project_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 tiny_user_project_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tiny_user_project_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tiny_user_project_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tiny_user_project_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tiny_user_project_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tiny_user_project_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tiny_user_project_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tiny_user_project_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tiny_user_project_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tiny_user_project_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tiny_user_project_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tiny_user_project_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 tiny_user_project_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 tiny_user_project_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 tiny_user_project_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 tiny_user_project_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 tiny_user_project_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 tiny_user_project_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 tiny_user_project_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 tiny_user_project_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 tiny_user_project_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 tiny_user_project_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 tiny_user_project_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 tiny_user_project_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 tiny_user_project_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 tiny_user_project_83 (.LO(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[10]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[10]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[8]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[9]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(io_out[21]));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(net3),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net2),
    .X(net13));
 sky130_fd_sc_hd__conb_1 tiny_user_project_14 (.LO(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[9]));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_297 ();
 assign io_oeb[0] = net14;
 assign io_oeb[10] = net24;
 assign io_oeb[11] = net25;
 assign io_oeb[12] = net26;
 assign io_oeb[13] = net27;
 assign io_oeb[14] = net28;
 assign io_oeb[15] = net29;
 assign io_oeb[16] = net30;
 assign io_oeb[17] = net31;
 assign io_oeb[18] = net32;
 assign io_oeb[19] = net33;
 assign io_oeb[1] = net15;
 assign io_oeb[20] = net34;
 assign io_oeb[21] = net35;
 assign io_oeb[22] = net36;
 assign io_oeb[23] = net37;
 assign io_oeb[24] = net38;
 assign io_oeb[25] = net39;
 assign io_oeb[26] = net40;
 assign io_oeb[27] = net41;
 assign io_oeb[28] = net42;
 assign io_oeb[29] = net43;
 assign io_oeb[2] = net16;
 assign io_oeb[30] = net44;
 assign io_oeb[31] = net45;
 assign io_oeb[32] = net46;
 assign io_oeb[33] = net47;
 assign io_oeb[34] = net48;
 assign io_oeb[35] = net49;
 assign io_oeb[36] = net50;
 assign io_oeb[37] = net51;
 assign io_oeb[3] = net17;
 assign io_oeb[4] = net18;
 assign io_oeb[5] = net19;
 assign io_oeb[6] = net20;
 assign io_oeb[7] = net21;
 assign io_oeb[8] = net22;
 assign io_oeb[9] = net23;
 assign io_out[0] = net52;
 assign io_out[10] = net62;
 assign io_out[11] = net63;
 assign io_out[12] = net64;
 assign io_out[13] = net65;
 assign io_out[14] = net66;
 assign io_out[15] = net67;
 assign io_out[1] = net53;
 assign io_out[22] = net68;
 assign io_out[23] = net69;
 assign io_out[24] = net70;
 assign io_out[25] = net71;
 assign io_out[26] = net72;
 assign io_out[27] = net73;
 assign io_out[28] = net74;
 assign io_out[29] = net75;
 assign io_out[2] = net54;
 assign io_out[30] = net76;
 assign io_out[31] = net77;
 assign io_out[32] = net78;
 assign io_out[33] = net79;
 assign io_out[34] = net80;
 assign io_out[35] = net81;
 assign io_out[36] = net82;
 assign io_out[37] = net83;
 assign io_out[3] = net55;
 assign io_out[4] = net56;
 assign io_out[5] = net57;
 assign io_out[6] = net58;
 assign io_out[7] = net59;
 assign io_out[8] = net60;
 assign io_out[9] = net61;
endmodule

