magic
tech sky130A
magscale 1 2
timestamp 1671710122
<< viali >>
rect 5089 17289 5123 17323
rect 5825 17289 5859 17323
rect 7665 17289 7699 17323
rect 17141 17221 17175 17255
rect 17601 17221 17635 17255
rect 2789 17153 2823 17187
rect 3433 17153 3467 17187
rect 5273 17153 5307 17187
rect 6009 17153 6043 17187
rect 6929 17153 6963 17187
rect 7481 17153 7515 17187
rect 8217 17153 8251 17187
rect 8585 17153 8619 17187
rect 9675 17153 9709 17187
rect 10425 17153 10459 17187
rect 10885 17153 10919 17187
rect 13737 17153 13771 17187
rect 16037 17153 16071 17187
rect 18337 17153 18371 17187
rect 8401 17085 8435 17119
rect 9597 17085 9631 17119
rect 11161 17085 11195 17119
rect 13461 17085 13495 17119
rect 15761 17085 15795 17119
rect 17049 17085 17083 17119
rect 4537 17017 4571 17051
rect 10701 17017 10735 17051
rect 17601 17017 17635 17051
rect 1593 16949 1627 16983
rect 6837 16949 6871 16983
rect 8309 16949 8343 16983
rect 8585 16949 8619 16983
rect 9873 16949 9907 16983
rect 10609 16949 10643 16983
rect 10793 16949 10827 16983
rect 11989 16949 12023 16983
rect 14289 16949 14323 16983
rect 16865 16949 16899 16983
rect 18153 16949 18187 16983
rect 2697 16745 2731 16779
rect 4721 16745 4755 16779
rect 10149 16745 10183 16779
rect 1593 16609 1627 16643
rect 10057 16609 10091 16643
rect 11069 16609 11103 16643
rect 11989 16609 12023 16643
rect 12265 16609 12299 16643
rect 14565 16609 14599 16643
rect 16773 16609 16807 16643
rect 5181 16541 5215 16575
rect 5365 16541 5399 16575
rect 7297 16541 7331 16575
rect 8033 16541 8067 16575
rect 8401 16541 8435 16575
rect 8585 16541 8619 16575
rect 9873 16541 9907 16575
rect 9965 16541 9999 16575
rect 10333 16541 10367 16575
rect 10793 16541 10827 16575
rect 10977 16541 11011 16575
rect 11161 16541 11195 16575
rect 11253 16541 11287 16575
rect 14289 16541 14323 16575
rect 16497 16541 16531 16575
rect 5273 16473 5307 16507
rect 6009 16473 6043 16507
rect 6653 16473 6687 16507
rect 6837 16473 6871 16507
rect 5917 16405 5951 16439
rect 7481 16405 7515 16439
rect 8401 16405 8435 16439
rect 9597 16405 9631 16439
rect 11529 16405 11563 16439
rect 13737 16405 13771 16439
rect 16037 16405 16071 16439
rect 18245 16405 18279 16439
rect 11161 16201 11195 16235
rect 16037 16201 16071 16235
rect 18153 16201 18187 16235
rect 6821 16133 6855 16167
rect 7021 16133 7055 16167
rect 13645 16133 13679 16167
rect 17049 16133 17083 16167
rect 17601 16133 17635 16167
rect 1593 16065 1627 16099
rect 2881 16065 2915 16099
rect 5181 16065 5215 16099
rect 5365 16065 5399 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 7573 16065 7607 16099
rect 7757 16065 7791 16099
rect 7941 16065 7975 16099
rect 8585 16065 8619 16099
rect 12541 16065 12575 16099
rect 13369 16065 13403 16099
rect 15853 16065 15887 16099
rect 18337 16065 18371 16099
rect 2237 15997 2271 16031
rect 8677 15997 8711 16031
rect 8953 15997 8987 16031
rect 9413 15997 9447 16031
rect 9689 15997 9723 16031
rect 12265 15997 12299 16031
rect 12449 15997 12483 16031
rect 15117 15997 15151 16031
rect 15945 15997 15979 16031
rect 16221 15997 16255 16031
rect 16313 15997 16347 16031
rect 17141 15997 17175 16031
rect 12909 15929 12943 15963
rect 15669 15929 15703 15963
rect 17601 15929 17635 15963
rect 5365 15861 5399 15895
rect 6009 15861 6043 15895
rect 6653 15861 6687 15895
rect 6837 15861 6871 15895
rect 7481 15861 7515 15895
rect 7665 15861 7699 15895
rect 16865 15861 16899 15895
rect 2237 15657 2271 15691
rect 6193 15657 6227 15691
rect 6653 15657 6687 15691
rect 9321 15657 9355 15691
rect 7573 15589 7607 15623
rect 8401 15589 8435 15623
rect 11529 15589 11563 15623
rect 11989 15589 12023 15623
rect 10057 15521 10091 15555
rect 13461 15521 13495 15555
rect 1593 15453 1627 15487
rect 6653 15453 6687 15487
rect 6837 15453 6871 15487
rect 7297 15453 7331 15487
rect 7573 15453 7607 15487
rect 8125 15453 8159 15487
rect 9781 15453 9815 15487
rect 13737 15453 13771 15487
rect 14335 15453 14369 15487
rect 15761 15453 15795 15487
rect 16129 15453 16163 15487
rect 16589 15453 16623 15487
rect 16865 15385 16899 15419
rect 8585 15317 8619 15351
rect 18337 15317 18371 15351
rect 7941 15113 7975 15147
rect 9045 15113 9079 15147
rect 12541 15113 12575 15147
rect 13001 15113 13035 15147
rect 8677 15045 8711 15079
rect 14473 15045 14507 15079
rect 15945 15045 15979 15079
rect 18061 15045 18095 15079
rect 1593 14977 1627 15011
rect 7205 14977 7239 15011
rect 7389 14977 7423 15011
rect 8125 14977 8159 15011
rect 8585 14977 8619 15011
rect 8861 14977 8895 15011
rect 9689 14977 9723 15011
rect 10517 14977 10551 15011
rect 10885 14977 10919 15011
rect 12173 14977 12207 15011
rect 14749 14977 14783 15011
rect 17417 14977 17451 15011
rect 18245 14977 18279 15011
rect 18337 14977 18371 15011
rect 9781 14909 9815 14943
rect 10057 14909 10091 14943
rect 10977 14909 11011 14943
rect 11897 14909 11931 14943
rect 12081 14909 12115 14943
rect 15393 14909 15427 14943
rect 15485 14909 15519 14943
rect 16865 14909 16899 14943
rect 17141 14909 17175 14943
rect 17509 14909 17543 14943
rect 7389 14841 7423 14875
rect 15945 14841 15979 14875
rect 6745 14773 6779 14807
rect 11161 14773 11195 14807
rect 15209 14773 15243 14807
rect 18061 14773 18095 14807
rect 7113 14569 7147 14603
rect 7941 14569 7975 14603
rect 8585 14569 8619 14603
rect 9413 14569 9447 14603
rect 11529 14569 11563 14603
rect 10149 14501 10183 14535
rect 10517 14501 10551 14535
rect 10057 14433 10091 14467
rect 11253 14433 11287 14467
rect 13737 14433 13771 14467
rect 14289 14433 14323 14467
rect 14565 14433 14599 14467
rect 16497 14433 16531 14467
rect 18245 14433 18279 14467
rect 1593 14365 1627 14399
rect 8401 14365 8435 14399
rect 10333 14365 10367 14399
rect 11161 14365 11195 14399
rect 9229 14297 9263 14331
rect 9445 14297 9479 14331
rect 13461 14297 13495 14331
rect 16773 14297 16807 14331
rect 9597 14229 9631 14263
rect 11989 14229 12023 14263
rect 16037 14229 16071 14263
rect 12909 14025 12943 14059
rect 16865 14025 16899 14059
rect 18127 14025 18161 14059
rect 9321 13957 9355 13991
rect 10977 13957 11011 13991
rect 12750 13957 12784 13991
rect 15945 13957 15979 13991
rect 16063 13957 16097 13991
rect 18337 13957 18371 13991
rect 8769 13889 8803 13923
rect 9229 13889 9263 13923
rect 9413 13889 9447 13923
rect 10057 13889 10091 13923
rect 10701 13889 10735 13923
rect 10885 13889 10919 13923
rect 11074 13889 11108 13923
rect 12253 13889 12287 13923
rect 12633 13889 12667 13923
rect 13369 13889 13403 13923
rect 15577 13889 15611 13923
rect 15761 13889 15795 13923
rect 15853 13889 15887 13923
rect 17049 13889 17083 13923
rect 17509 13889 17543 13923
rect 1593 13821 1627 13855
rect 9873 13821 9907 13855
rect 12541 13821 12575 13855
rect 13645 13821 13679 13855
rect 16221 13821 16255 13855
rect 17141 13821 17175 13855
rect 10241 13685 10275 13719
rect 10701 13685 10735 13719
rect 15117 13685 15151 13719
rect 17417 13685 17451 13719
rect 17969 13685 18003 13719
rect 18153 13685 18187 13719
rect 9965 13481 9999 13515
rect 12265 13481 12299 13515
rect 17049 13481 17083 13515
rect 17601 13481 17635 13515
rect 17877 13481 17911 13515
rect 10609 13413 10643 13447
rect 11345 13345 11379 13379
rect 13093 13345 13127 13379
rect 13369 13345 13403 13379
rect 17877 13345 17911 13379
rect 1593 13277 1627 13311
rect 9781 13277 9815 13311
rect 9965 13277 9999 13311
rect 10425 13277 10459 13311
rect 10517 13277 10551 13311
rect 10701 13277 10735 13311
rect 11161 13277 11195 13311
rect 11483 13277 11517 13311
rect 11621 13277 11655 13311
rect 12633 13277 12667 13311
rect 13277 13277 13311 13311
rect 14289 13277 14323 13311
rect 16681 13277 16715 13311
rect 16773 13277 16807 13311
rect 18153 13277 18187 13311
rect 12265 13209 12299 13243
rect 14565 13209 14599 13243
rect 17141 13209 17175 13243
rect 11253 13141 11287 13175
rect 12081 13141 12115 13175
rect 13737 13141 13771 13175
rect 16037 13141 16071 13175
rect 16497 13141 16531 13175
rect 12265 12937 12299 12971
rect 17417 12937 17451 12971
rect 14013 12869 14047 12903
rect 16097 12869 16131 12903
rect 16313 12869 16347 12903
rect 10517 12801 10551 12835
rect 10977 12801 11011 12835
rect 11161 12801 11195 12835
rect 11805 12801 11839 12835
rect 12081 12801 12115 12835
rect 12909 12801 12943 12835
rect 16865 12801 16899 12835
rect 17233 12801 17267 12835
rect 17877 12801 17911 12835
rect 12817 12733 12851 12767
rect 13277 12733 13311 12767
rect 13737 12733 13771 12767
rect 17969 12733 18003 12767
rect 10977 12665 11011 12699
rect 15945 12665 15979 12699
rect 18245 12665 18279 12699
rect 1593 12597 1627 12631
rect 11897 12597 11931 12631
rect 15485 12597 15519 12631
rect 16129 12597 16163 12631
rect 17233 12597 17267 12631
rect 17969 12597 18003 12631
rect 12357 12393 12391 12427
rect 15025 12393 15059 12427
rect 16773 12393 16807 12427
rect 13737 12325 13771 12359
rect 15761 12325 15795 12359
rect 16865 12325 16899 12359
rect 17785 12325 17819 12359
rect 12725 12257 12759 12291
rect 1593 12189 1627 12223
rect 11805 12189 11839 12223
rect 11897 12189 11931 12223
rect 12541 12189 12575 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 13553 12189 13587 12223
rect 14657 12189 14691 12223
rect 15025 12189 15059 12223
rect 15301 12189 15335 12223
rect 15945 12189 15979 12223
rect 16037 12189 16071 12223
rect 16313 12189 16347 12223
rect 17969 12189 18003 12223
rect 13461 12121 13495 12155
rect 14815 12121 14849 12155
rect 16129 12121 16163 12155
rect 17233 12121 17267 12155
rect 13093 11849 13127 11883
rect 13921 11849 13955 11883
rect 18153 11849 18187 11883
rect 14197 11781 14231 11815
rect 17141 11781 17175 11815
rect 12633 11713 12667 11747
rect 13277 11713 13311 11747
rect 14105 11713 14139 11747
rect 14289 11713 14323 11747
rect 14473 11713 14507 11747
rect 15117 11713 15151 11747
rect 15485 11713 15519 11747
rect 15945 11713 15979 11747
rect 16037 11713 16071 11747
rect 16957 11713 16991 11747
rect 17693 11713 17727 11747
rect 18337 11713 18371 11747
rect 13461 11645 13495 11679
rect 1593 11509 1627 11543
rect 14933 11509 14967 11543
rect 15393 11509 15427 11543
rect 15945 11509 15979 11543
rect 16313 11509 16347 11543
rect 13645 11305 13679 11339
rect 14289 11305 14323 11339
rect 15301 11305 15335 11339
rect 16313 11305 16347 11339
rect 17141 11305 17175 11339
rect 18337 11305 18371 11339
rect 14473 11237 14507 11271
rect 14749 11169 14783 11203
rect 16129 11169 16163 11203
rect 13553 11101 13587 11135
rect 13737 11101 13771 11135
rect 16221 11101 16255 11135
rect 16957 11101 16991 11135
rect 15577 11033 15611 11067
rect 16497 11033 16531 11067
rect 16405 10965 16439 10999
rect 14197 10761 14231 10795
rect 15117 10761 15151 10795
rect 15577 10761 15611 10795
rect 16957 10761 16991 10795
rect 14289 10625 14323 10659
rect 14749 10625 14783 10659
rect 15853 10625 15887 10659
rect 15945 10625 15979 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 17693 10625 17727 10659
rect 18337 10625 18371 10659
rect 1593 10557 1627 10591
rect 14841 10557 14875 10591
rect 14933 10421 14967 10455
rect 15945 10421 15979 10455
rect 15945 10217 15979 10251
rect 17049 10217 17083 10251
rect 17509 10217 17543 10251
rect 18337 10217 18371 10251
rect 1593 10149 1627 10183
rect 15117 10149 15151 10183
rect 14933 10013 14967 10047
rect 15117 10013 15151 10047
rect 17693 10013 17727 10047
rect 16313 9537 16347 9571
rect 17693 9537 17727 9571
rect 18337 9537 18371 9571
rect 15669 9469 15703 9503
rect 17049 9469 17083 9503
rect 18153 9401 18187 9435
rect 1593 9333 1627 9367
rect 17693 9129 17727 9163
rect 18337 9129 18371 9163
rect 16405 9061 16439 9095
rect 1593 8925 1627 8959
rect 17049 8925 17083 8959
rect 17049 8449 17083 8483
rect 17693 8449 17727 8483
rect 18337 8449 18371 8483
rect 1593 8313 1627 8347
rect 17693 8041 17727 8075
rect 18337 7905 18371 7939
rect 1593 7837 1627 7871
rect 18337 7361 18371 7395
rect 1593 7157 1627 7191
rect 1593 6749 1627 6783
rect 18337 6749 18371 6783
rect 18337 6273 18371 6307
rect 1593 5661 1627 5695
rect 18337 5661 18371 5695
rect 1593 5185 1627 5219
rect 18337 5049 18371 5083
rect 1593 4573 1627 4607
rect 18337 4573 18371 4607
rect 1593 4029 1627 4063
rect 18337 3893 18371 3927
rect 1593 3485 1627 3519
rect 18337 3485 18371 3519
rect 1593 2805 1627 2839
rect 18337 2805 18371 2839
rect 1593 2397 1627 2431
rect 2237 2397 2271 2431
rect 17693 2397 17727 2431
rect 18337 2397 18371 2431
<< metal1 >>
rect 8110 17824 8116 17876
rect 8168 17864 8174 17876
rect 10410 17864 10416 17876
rect 8168 17836 10416 17864
rect 8168 17824 8174 17836
rect 10410 17824 10416 17836
rect 10468 17864 10474 17876
rect 17126 17864 17132 17876
rect 10468 17836 17132 17864
rect 10468 17824 10474 17836
rect 17126 17824 17132 17836
rect 17184 17824 17190 17876
rect 6178 17756 6184 17808
rect 6236 17796 6242 17808
rect 14642 17796 14648 17808
rect 6236 17768 14648 17796
rect 6236 17756 6242 17768
rect 14642 17756 14648 17768
rect 14700 17756 14706 17808
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 13722 17728 13728 17740
rect 9456 17700 13728 17728
rect 9456 17688 9462 17700
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 8478 17552 8484 17604
rect 8536 17592 8542 17604
rect 10226 17592 10232 17604
rect 8536 17564 10232 17592
rect 8536 17552 8542 17564
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 4706 17484 4712 17536
rect 4764 17524 4770 17536
rect 13630 17524 13636 17536
rect 4764 17496 13636 17524
rect 4764 17484 4770 17496
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 1104 17434 19019 17456
rect 1104 17382 5388 17434
rect 5440 17382 5452 17434
rect 5504 17382 5516 17434
rect 5568 17382 5580 17434
rect 5632 17382 5644 17434
rect 5696 17382 9827 17434
rect 9879 17382 9891 17434
rect 9943 17382 9955 17434
rect 10007 17382 10019 17434
rect 10071 17382 10083 17434
rect 10135 17382 14266 17434
rect 14318 17382 14330 17434
rect 14382 17382 14394 17434
rect 14446 17382 14458 17434
rect 14510 17382 14522 17434
rect 14574 17382 18705 17434
rect 18757 17382 18769 17434
rect 18821 17382 18833 17434
rect 18885 17382 18897 17434
rect 18949 17382 18961 17434
rect 19013 17382 19019 17434
rect 1104 17360 19019 17382
rect 5077 17323 5135 17329
rect 5077 17289 5089 17323
rect 5123 17320 5135 17323
rect 5718 17320 5724 17332
rect 5123 17292 5724 17320
rect 5123 17289 5135 17292
rect 5077 17283 5135 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 7558 17320 7564 17332
rect 5859 17292 7564 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17320 7711 17323
rect 11790 17320 11796 17332
rect 7699 17292 11796 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 14182 17320 14188 17332
rect 11900 17292 14188 17320
rect 8110 17212 8116 17264
rect 8168 17212 8174 17264
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 11900 17252 11928 17292
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 14274 17280 14280 17332
rect 14332 17320 14338 17332
rect 14332 17292 16068 17320
rect 14332 17280 14338 17292
rect 8352 17224 11928 17252
rect 8352 17212 8358 17224
rect 12986 17212 12992 17264
rect 13044 17212 13050 17264
rect 14734 17212 14740 17264
rect 14792 17212 14798 17264
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 3326 17184 3332 17196
rect 2823 17156 3332 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17184 3479 17187
rect 4798 17184 4804 17196
rect 3467 17156 4804 17184
rect 3467 17153 3479 17156
rect 3421 17147 3479 17153
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 5166 17144 5172 17196
rect 5224 17184 5230 17196
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 5224 17156 5273 17184
rect 5224 17144 5230 17156
rect 5261 17153 5273 17156
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17153 6055 17187
rect 6914 17184 6920 17196
rect 6875 17156 6920 17184
rect 5997 17147 6055 17153
rect 6012 17116 6040 17147
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 7469 17187 7527 17193
rect 7469 17184 7481 17187
rect 7432 17156 7481 17184
rect 7432 17144 7438 17156
rect 7469 17153 7481 17156
rect 7515 17153 7527 17187
rect 8128 17184 8156 17212
rect 8205 17187 8263 17193
rect 8205 17184 8217 17187
rect 8128 17156 8217 17184
rect 7469 17147 7527 17153
rect 8205 17153 8217 17156
rect 8251 17153 8263 17187
rect 8570 17184 8576 17196
rect 8531 17156 8576 17184
rect 8205 17147 8263 17153
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 9663 17187 9721 17193
rect 9663 17153 9675 17187
rect 9709 17153 9721 17187
rect 10410 17184 10416 17196
rect 10371 17156 10416 17184
rect 9663 17147 9721 17153
rect 8386 17116 8392 17128
rect 6012 17088 8392 17116
rect 8386 17076 8392 17088
rect 8444 17116 8450 17128
rect 9585 17119 9643 17125
rect 8444 17088 8537 17116
rect 8444 17076 8450 17088
rect 9585 17085 9597 17119
rect 9631 17085 9643 17119
rect 9692 17116 9720 17147
rect 10410 17144 10416 17156
rect 10468 17144 10474 17196
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 10520 17156 10885 17184
rect 10520 17116 10548 17156
rect 10873 17153 10885 17156
rect 10919 17184 10931 17187
rect 11054 17184 11060 17196
rect 10919 17156 11060 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 16040 17193 16068 17292
rect 17034 17212 17040 17264
rect 17092 17252 17098 17264
rect 17129 17255 17187 17261
rect 17129 17252 17141 17255
rect 17092 17224 17141 17252
rect 17092 17212 17098 17224
rect 17129 17221 17141 17224
rect 17175 17221 17187 17255
rect 17129 17215 17187 17221
rect 17218 17212 17224 17264
rect 17276 17252 17282 17264
rect 17589 17255 17647 17261
rect 17589 17252 17601 17255
rect 17276 17224 17601 17252
rect 17276 17212 17282 17224
rect 17589 17221 17601 17224
rect 17635 17221 17647 17255
rect 17589 17215 17647 17221
rect 16025 17187 16083 17193
rect 13780 17156 13825 17184
rect 13780 17144 13786 17156
rect 16025 17153 16037 17187
rect 16071 17153 16083 17187
rect 18322 17184 18328 17196
rect 18283 17156 18328 17184
rect 16025 17147 16083 17153
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 9692 17088 10548 17116
rect 11149 17119 11207 17125
rect 9585 17079 9643 17085
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 12802 17116 12808 17128
rect 11195 17088 12808 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 4525 17051 4583 17057
rect 4525 17017 4537 17051
rect 4571 17048 4583 17051
rect 9214 17048 9220 17060
rect 4571 17020 9220 17048
rect 4571 17017 4583 17020
rect 4525 17011 4583 17017
rect 9214 17008 9220 17020
rect 9272 17008 9278 17060
rect 9600 17048 9628 17079
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 13446 17116 13452 17128
rect 13407 17088 13452 17116
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 14182 17076 14188 17128
rect 14240 17116 14246 17128
rect 15749 17119 15807 17125
rect 15749 17116 15761 17119
rect 14240 17088 15761 17116
rect 14240 17076 14246 17088
rect 15749 17085 15761 17088
rect 15795 17085 15807 17119
rect 15749 17079 15807 17085
rect 16390 17076 16396 17128
rect 16448 17116 16454 17128
rect 17037 17119 17095 17125
rect 17037 17116 17049 17119
rect 16448 17088 17049 17116
rect 16448 17076 16454 17088
rect 17037 17085 17049 17088
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 9416 17020 9628 17048
rect 10689 17051 10747 17057
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 1452 16952 1593 16980
rect 1452 16940 1458 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 6825 16983 6883 16989
rect 6825 16980 6837 16983
rect 6696 16952 6837 16980
rect 6696 16940 6702 16952
rect 6825 16949 6837 16952
rect 6871 16949 6883 16983
rect 6825 16943 6883 16949
rect 7098 16940 7104 16992
rect 7156 16980 7162 16992
rect 8297 16983 8355 16989
rect 8297 16980 8309 16983
rect 7156 16952 8309 16980
rect 7156 16940 7162 16952
rect 8297 16949 8309 16952
rect 8343 16980 8355 16983
rect 8478 16980 8484 16992
rect 8343 16952 8484 16980
rect 8343 16949 8355 16952
rect 8297 16943 8355 16949
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 8573 16983 8631 16989
rect 8573 16949 8585 16983
rect 8619 16980 8631 16983
rect 9122 16980 9128 16992
rect 8619 16952 9128 16980
rect 8619 16949 8631 16952
rect 8573 16943 8631 16949
rect 9122 16940 9128 16952
rect 9180 16980 9186 16992
rect 9416 16980 9444 17020
rect 10689 17017 10701 17051
rect 10735 17048 10747 17051
rect 11054 17048 11060 17060
rect 10735 17020 11060 17048
rect 10735 17017 10747 17020
rect 10689 17011 10747 17017
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 17586 17048 17592 17060
rect 15948 17020 16988 17048
rect 17547 17020 17592 17048
rect 9180 16952 9444 16980
rect 9180 16940 9186 16952
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 9861 16983 9919 16989
rect 9861 16980 9873 16983
rect 9732 16952 9873 16980
rect 9732 16940 9738 16952
rect 9861 16949 9873 16952
rect 9907 16949 9919 16983
rect 9861 16943 9919 16949
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10597 16983 10655 16989
rect 10597 16980 10609 16983
rect 10284 16952 10609 16980
rect 10284 16940 10290 16952
rect 10597 16949 10609 16952
rect 10643 16949 10655 16983
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10597 16943 10655 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 10870 16940 10876 16992
rect 10928 16980 10934 16992
rect 11977 16983 12035 16989
rect 11977 16980 11989 16983
rect 10928 16952 11989 16980
rect 10928 16940 10934 16952
rect 11977 16949 11989 16952
rect 12023 16949 12035 16983
rect 11977 16943 12035 16949
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 14277 16983 14335 16989
rect 14277 16980 14289 16983
rect 13780 16952 14289 16980
rect 13780 16940 13786 16952
rect 14277 16949 14289 16952
rect 14323 16949 14335 16983
rect 14277 16943 14335 16949
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 15948 16980 15976 17020
rect 16850 16980 16856 16992
rect 14700 16952 15976 16980
rect 16811 16952 16856 16980
rect 14700 16940 14706 16952
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 16960 16980 16988 17020
rect 17586 17008 17592 17020
rect 17644 17008 17650 17060
rect 18141 16983 18199 16989
rect 18141 16980 18153 16983
rect 16960 16952 18153 16980
rect 18141 16949 18153 16952
rect 18187 16949 18199 16983
rect 18141 16943 18199 16949
rect 1104 16890 18860 16912
rect 1104 16838 3169 16890
rect 3221 16838 3233 16890
rect 3285 16838 3297 16890
rect 3349 16838 3361 16890
rect 3413 16838 3425 16890
rect 3477 16838 7608 16890
rect 7660 16838 7672 16890
rect 7724 16838 7736 16890
rect 7788 16838 7800 16890
rect 7852 16838 7864 16890
rect 7916 16838 12047 16890
rect 12099 16838 12111 16890
rect 12163 16838 12175 16890
rect 12227 16838 12239 16890
rect 12291 16838 12303 16890
rect 12355 16838 16486 16890
rect 16538 16838 16550 16890
rect 16602 16838 16614 16890
rect 16666 16838 16678 16890
rect 16730 16838 16742 16890
rect 16794 16838 18860 16890
rect 1104 16816 18860 16838
rect 2590 16736 2596 16788
rect 2648 16776 2654 16788
rect 2685 16779 2743 16785
rect 2685 16776 2697 16779
rect 2648 16748 2697 16776
rect 2648 16736 2654 16748
rect 2685 16745 2697 16748
rect 2731 16745 2743 16779
rect 4706 16776 4712 16788
rect 4667 16748 4712 16776
rect 2685 16739 2743 16745
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 8110 16776 8116 16788
rect 5920 16748 8116 16776
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 5920 16640 5948 16748
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 8386 16736 8392 16788
rect 8444 16776 8450 16788
rect 10042 16776 10048 16788
rect 8444 16748 10048 16776
rect 8444 16736 8450 16748
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 10226 16776 10232 16788
rect 10183 16748 10232 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 10226 16736 10232 16748
rect 10284 16736 10290 16788
rect 10318 16736 10324 16788
rect 10376 16776 10382 16788
rect 13446 16776 13452 16788
rect 10376 16748 13452 16776
rect 10376 16736 10382 16748
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 13906 16736 13912 16788
rect 13964 16776 13970 16788
rect 16114 16776 16120 16788
rect 13964 16748 16120 16776
rect 13964 16736 13970 16748
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 6638 16668 6644 16720
rect 6696 16708 6702 16720
rect 6696 16680 12020 16708
rect 6696 16668 6702 16680
rect 5736 16612 5948 16640
rect 8496 16612 8708 16640
rect 5166 16572 5172 16584
rect 5079 16544 5172 16572
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5353 16575 5411 16581
rect 5353 16541 5365 16575
rect 5399 16572 5411 16575
rect 5736 16572 5764 16612
rect 7285 16575 7343 16581
rect 7285 16572 7297 16575
rect 5399 16544 5764 16572
rect 5828 16544 7297 16572
rect 5399 16541 5411 16544
rect 5353 16535 5411 16541
rect 5184 16436 5212 16532
rect 5261 16507 5319 16513
rect 5261 16473 5273 16507
rect 5307 16504 5319 16507
rect 5828 16504 5856 16544
rect 7285 16541 7297 16544
rect 7331 16541 7343 16575
rect 8018 16572 8024 16584
rect 7979 16544 8024 16572
rect 7285 16535 7343 16541
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 8294 16532 8300 16584
rect 8352 16572 8358 16584
rect 8389 16575 8447 16581
rect 8389 16572 8401 16575
rect 8352 16544 8401 16572
rect 8352 16532 8358 16544
rect 8389 16541 8401 16544
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 5994 16504 6000 16516
rect 5307 16476 5856 16504
rect 5955 16476 6000 16504
rect 5307 16473 5319 16476
rect 5261 16467 5319 16473
rect 5994 16464 6000 16476
rect 6052 16464 6058 16516
rect 6638 16504 6644 16516
rect 6599 16476 6644 16504
rect 6638 16464 6644 16476
rect 6696 16464 6702 16516
rect 6825 16507 6883 16513
rect 6825 16473 6837 16507
rect 6871 16504 6883 16507
rect 7834 16504 7840 16516
rect 6871 16476 7840 16504
rect 6871 16473 6883 16476
rect 6825 16467 6883 16473
rect 7834 16464 7840 16476
rect 7892 16464 7898 16516
rect 8496 16504 8524 16612
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16541 8631 16575
rect 8573 16535 8631 16541
rect 8266 16476 8524 16504
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 5184 16408 5917 16436
rect 5905 16405 5917 16408
rect 5951 16436 5963 16439
rect 7098 16436 7104 16448
rect 5951 16408 7104 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 7469 16439 7527 16445
rect 7469 16405 7481 16439
rect 7515 16436 7527 16439
rect 8266 16436 8294 16476
rect 8386 16436 8392 16448
rect 7515 16408 8294 16436
rect 8347 16408 8392 16436
rect 7515 16405 7527 16408
rect 7469 16399 7527 16405
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 8588 16436 8616 16535
rect 8680 16504 8708 16612
rect 8754 16600 8760 16652
rect 8812 16640 8818 16652
rect 8812 16612 9996 16640
rect 8812 16600 8818 16612
rect 9968 16581 9996 16612
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 11054 16640 11060 16652
rect 10100 16612 11060 16640
rect 10100 16600 10106 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 11992 16649 12020 16680
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16609 12035 16643
rect 12250 16640 12256 16652
rect 12211 16612 12256 16640
rect 11977 16603 12035 16609
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 9953 16575 10011 16581
rect 9953 16541 9965 16575
rect 9999 16541 10011 16575
rect 9953 16535 10011 16541
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 10410 16572 10416 16584
rect 10367 16544 10416 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 9766 16504 9772 16516
rect 8680 16476 9772 16504
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 9306 16436 9312 16448
rect 8588 16408 9312 16436
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9582 16436 9588 16448
rect 9543 16408 9588 16436
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 9876 16436 9904 16535
rect 9968 16504 9996 16535
rect 10410 16532 10416 16544
rect 10468 16572 10474 16584
rect 10781 16575 10839 16581
rect 10781 16572 10793 16575
rect 10468 16544 10793 16572
rect 10468 16532 10474 16544
rect 10781 16541 10793 16544
rect 10827 16541 10839 16575
rect 10962 16572 10968 16584
rect 10923 16544 10968 16572
rect 10781 16535 10839 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11149 16575 11207 16581
rect 11149 16541 11161 16575
rect 11195 16541 11207 16575
rect 11149 16535 11207 16541
rect 11241 16575 11299 16581
rect 11241 16541 11253 16575
rect 11287 16572 11299 16575
rect 11330 16572 11336 16584
rect 11287 16544 11336 16572
rect 11287 16541 11299 16544
rect 11241 16535 11299 16541
rect 10594 16504 10600 16516
rect 9968 16476 10600 16504
rect 10594 16464 10600 16476
rect 10652 16504 10658 16516
rect 11164 16504 11192 16535
rect 11330 16532 11336 16544
rect 11388 16532 11394 16584
rect 10652 16476 11192 16504
rect 10652 16464 10658 16476
rect 10686 16436 10692 16448
rect 9876 16408 10692 16436
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 11517 16439 11575 16445
rect 11517 16405 11529 16439
rect 11563 16436 11575 16439
rect 11882 16436 11888 16448
rect 11563 16408 11888 16436
rect 11563 16405 11575 16408
rect 11517 16399 11575 16405
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 11992 16436 12020 16603
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 12400 16612 14565 16640
rect 12400 16600 12406 16612
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 14918 16600 14924 16652
rect 14976 16640 14982 16652
rect 16758 16640 16764 16652
rect 14976 16612 15792 16640
rect 16719 16612 16764 16640
rect 14976 16600 14982 16612
rect 13538 16532 13544 16584
rect 13596 16572 13602 16584
rect 14274 16572 14280 16584
rect 13596 16544 14280 16572
rect 13596 16532 13602 16544
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 15764 16572 15792 16612
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 15764 16544 15884 16572
rect 13998 16504 14004 16516
rect 13478 16476 14004 16504
rect 13998 16464 14004 16476
rect 14056 16504 14062 16516
rect 15856 16504 15884 16544
rect 16114 16532 16120 16584
rect 16172 16572 16178 16584
rect 16485 16575 16543 16581
rect 16485 16572 16497 16575
rect 16172 16544 16497 16572
rect 16172 16532 16178 16544
rect 16485 16541 16497 16544
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 14056 16476 15042 16504
rect 15856 16476 16160 16504
rect 14056 16464 14062 16476
rect 14752 16448 14780 16476
rect 13170 16436 13176 16448
rect 11992 16408 13176 16436
rect 13170 16396 13176 16408
rect 13228 16436 13234 16448
rect 13538 16436 13544 16448
rect 13228 16408 13544 16436
rect 13228 16396 13234 16408
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 13725 16439 13783 16445
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 13814 16436 13820 16448
rect 13771 16408 13820 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 14734 16396 14740 16448
rect 14792 16396 14798 16448
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 16025 16439 16083 16445
rect 16025 16436 16037 16439
rect 15528 16408 16037 16436
rect 15528 16396 15534 16408
rect 16025 16405 16037 16408
rect 16071 16405 16083 16439
rect 16132 16436 16160 16476
rect 17310 16464 17316 16516
rect 17368 16464 17374 16516
rect 18322 16504 18328 16516
rect 18064 16476 18328 16504
rect 18064 16436 18092 16476
rect 18322 16464 18328 16476
rect 18380 16464 18386 16516
rect 18230 16436 18236 16448
rect 16132 16408 18092 16436
rect 18191 16408 18236 16436
rect 16025 16399 16083 16405
rect 18230 16396 18236 16408
rect 18288 16396 18294 16448
rect 1104 16346 19019 16368
rect 1104 16294 5388 16346
rect 5440 16294 5452 16346
rect 5504 16294 5516 16346
rect 5568 16294 5580 16346
rect 5632 16294 5644 16346
rect 5696 16294 9827 16346
rect 9879 16294 9891 16346
rect 9943 16294 9955 16346
rect 10007 16294 10019 16346
rect 10071 16294 10083 16346
rect 10135 16294 14266 16346
rect 14318 16294 14330 16346
rect 14382 16294 14394 16346
rect 14446 16294 14458 16346
rect 14510 16294 14522 16346
rect 14574 16294 18705 16346
rect 18757 16294 18769 16346
rect 18821 16294 18833 16346
rect 18885 16294 18897 16346
rect 18949 16294 18961 16346
rect 19013 16294 19019 16346
rect 1104 16272 19019 16294
rect 5828 16204 8524 16232
rect 1118 16056 1124 16108
rect 1176 16096 1182 16108
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 1176 16068 1593 16096
rect 1176 16056 1182 16068
rect 1581 16065 1593 16068
rect 1627 16065 1639 16099
rect 2866 16096 2872 16108
rect 2827 16068 2872 16096
rect 1581 16059 1639 16065
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 5166 16096 5172 16108
rect 5127 16068 5172 16096
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 5350 16096 5356 16108
rect 5311 16068 5356 16096
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 5828 16105 5856 16204
rect 6822 16173 6828 16176
rect 6809 16167 6828 16173
rect 6809 16133 6821 16167
rect 6809 16127 6828 16133
rect 6822 16124 6828 16127
rect 6880 16124 6886 16176
rect 7009 16167 7067 16173
rect 7009 16133 7021 16167
rect 7055 16164 7067 16167
rect 7098 16164 7104 16176
rect 7055 16136 7104 16164
rect 7055 16133 7067 16136
rect 7009 16127 7067 16133
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 7190 16124 7196 16176
rect 7248 16164 7254 16176
rect 8496 16164 8524 16204
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 11149 16235 11207 16241
rect 8628 16204 11100 16232
rect 8628 16192 8634 16204
rect 9950 16164 9956 16176
rect 7248 16136 8432 16164
rect 8496 16136 9956 16164
rect 7248 16124 7254 16136
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5997 16099 6055 16105
rect 5997 16065 6009 16099
rect 6043 16065 6055 16099
rect 7561 16099 7619 16105
rect 7561 16096 7573 16099
rect 5997 16059 6055 16065
rect 7484 16068 7573 16096
rect 382 15988 388 16040
rect 440 16028 446 16040
rect 2225 16031 2283 16037
rect 2225 16028 2237 16031
rect 440 16000 2237 16028
rect 440 15988 446 16000
rect 2225 15997 2237 16000
rect 2271 15997 2283 16031
rect 2225 15991 2283 15997
rect 6012 15960 6040 16059
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 7484 16028 7512 16068
rect 7561 16065 7573 16068
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 7929 16099 7987 16105
rect 7800 16068 7845 16096
rect 7800 16056 7806 16068
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 8294 16096 8300 16108
rect 7975 16068 8300 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8404 16096 8432 16136
rect 9950 16124 9956 16136
rect 10008 16124 10014 16176
rect 11072 16164 11100 16204
rect 11149 16201 11161 16235
rect 11195 16232 11207 16235
rect 13262 16232 13268 16244
rect 11195 16204 13268 16232
rect 11195 16201 11207 16204
rect 11149 16195 11207 16201
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 15838 16232 15844 16244
rect 13872 16204 15844 16232
rect 13872 16192 13878 16204
rect 15838 16192 15844 16204
rect 15896 16232 15902 16244
rect 16025 16235 16083 16241
rect 16025 16232 16037 16235
rect 15896 16204 16037 16232
rect 15896 16192 15902 16204
rect 16025 16201 16037 16204
rect 16071 16201 16083 16235
rect 18141 16235 18199 16241
rect 18141 16232 18153 16235
rect 16025 16195 16083 16201
rect 16132 16204 18153 16232
rect 13633 16167 13691 16173
rect 13633 16164 13645 16167
rect 11072 16136 13645 16164
rect 13633 16133 13645 16136
rect 13679 16133 13691 16167
rect 13633 16127 13691 16133
rect 14918 16124 14924 16176
rect 14976 16164 14982 16176
rect 16132 16164 16160 16204
rect 18141 16201 18153 16204
rect 18187 16201 18199 16235
rect 18141 16195 18199 16201
rect 17034 16164 17040 16176
rect 14976 16136 16160 16164
rect 16995 16136 17040 16164
rect 14976 16124 14982 16136
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 17586 16164 17592 16176
rect 17547 16136 17592 16164
rect 17586 16124 17592 16136
rect 17644 16124 17650 16176
rect 8573 16099 8631 16105
rect 8573 16096 8585 16099
rect 8404 16068 8585 16096
rect 8573 16065 8585 16068
rect 8619 16096 8631 16099
rect 9030 16096 9036 16108
rect 8619 16068 9036 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 10778 16056 10784 16108
rect 10836 16056 10842 16108
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 11020 16068 11376 16096
rect 11020 16056 11026 16068
rect 6696 16000 7512 16028
rect 6696 15988 6702 16000
rect 7834 15988 7840 16040
rect 7892 16028 7898 16040
rect 7892 16000 8616 16028
rect 7892 15988 7898 16000
rect 8588 15960 8616 16000
rect 8662 15988 8668 16040
rect 8720 16028 8726 16040
rect 8938 16028 8944 16040
rect 8720 16000 8765 16028
rect 8899 16000 8944 16028
rect 8720 15988 8726 16000
rect 8938 15988 8944 16000
rect 8996 15988 9002 16040
rect 9398 16028 9404 16040
rect 9048 16000 9404 16028
rect 9048 15960 9076 16000
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 9723 16000 11284 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 6012 15932 8340 15960
rect 8588 15932 9076 15960
rect 5258 15852 5264 15904
rect 5316 15892 5322 15904
rect 5353 15895 5411 15901
rect 5353 15892 5365 15895
rect 5316 15864 5365 15892
rect 5316 15852 5322 15864
rect 5353 15861 5365 15864
rect 5399 15861 5411 15895
rect 5994 15892 6000 15904
rect 5955 15864 6000 15892
rect 5353 15855 5411 15861
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 6730 15892 6736 15904
rect 6687 15864 6736 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 7466 15892 7472 15904
rect 6880 15864 6925 15892
rect 7427 15864 7472 15892
rect 6880 15852 6886 15864
rect 7466 15852 7472 15864
rect 7524 15852 7530 15904
rect 7653 15895 7711 15901
rect 7653 15861 7665 15895
rect 7699 15892 7711 15895
rect 8202 15892 8208 15904
rect 7699 15864 8208 15892
rect 7699 15861 7711 15864
rect 7653 15855 7711 15861
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 8312 15892 8340 15932
rect 10410 15892 10416 15904
rect 8312 15864 10416 15892
rect 10410 15852 10416 15864
rect 10468 15892 10474 15904
rect 10870 15892 10876 15904
rect 10468 15864 10876 15892
rect 10468 15852 10474 15864
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 11256 15892 11284 16000
rect 11348 15960 11376 16068
rect 11790 16056 11796 16108
rect 11848 16096 11854 16108
rect 12529 16099 12587 16105
rect 12529 16096 12541 16099
rect 11848 16068 12541 16096
rect 11848 16056 11854 16068
rect 12529 16065 12541 16068
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 13228 16068 13369 16096
rect 13228 16056 13234 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 14734 16056 14740 16108
rect 14792 16056 14798 16108
rect 15838 16096 15844 16108
rect 15799 16068 15844 16096
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 18325 16099 18383 16105
rect 18325 16096 18337 16099
rect 16040 16068 18337 16096
rect 11882 15988 11888 16040
rect 11940 16028 11946 16040
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 11940 16000 12265 16028
rect 11940 15988 11946 16000
rect 12253 15997 12265 16000
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 14826 16028 14832 16040
rect 12437 15991 12495 15997
rect 13464 16000 14832 16028
rect 12452 15960 12480 15991
rect 11348 15932 12480 15960
rect 12897 15963 12955 15969
rect 12897 15929 12909 15963
rect 12943 15960 12955 15963
rect 13464 15960 13492 16000
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15010 15988 15016 16040
rect 15068 16028 15074 16040
rect 15105 16031 15163 16037
rect 15105 16028 15117 16031
rect 15068 16000 15117 16028
rect 15068 15988 15074 16000
rect 15105 15997 15117 16000
rect 15151 15997 15163 16031
rect 15105 15991 15163 15997
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 15933 16031 15991 16037
rect 15933 16028 15945 16031
rect 15436 16000 15945 16028
rect 15436 15988 15442 16000
rect 15933 15997 15945 16000
rect 15979 15997 15991 16031
rect 15933 15991 15991 15997
rect 12943 15932 13492 15960
rect 12943 15929 12955 15932
rect 12897 15923 12955 15929
rect 14642 15920 14648 15972
rect 14700 15960 14706 15972
rect 15657 15963 15715 15969
rect 15657 15960 15669 15963
rect 14700 15932 15669 15960
rect 14700 15920 14706 15932
rect 15657 15929 15669 15932
rect 15703 15929 15715 15963
rect 15657 15923 15715 15929
rect 12434 15892 12440 15904
rect 11256 15864 12440 15892
rect 12434 15852 12440 15864
rect 12492 15852 12498 15904
rect 12526 15852 12532 15904
rect 12584 15892 12590 15904
rect 16040 15892 16068 16068
rect 18325 16065 18337 16068
rect 18371 16065 18383 16099
rect 18325 16059 18383 16065
rect 16206 16028 16212 16040
rect 16167 16000 16212 16028
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 17129 16031 17187 16037
rect 16356 16000 16401 16028
rect 16356 15988 16362 16000
rect 17129 15997 17141 16031
rect 17175 16028 17187 16031
rect 17218 16028 17224 16040
rect 17175 16000 17224 16028
rect 17175 15997 17187 16000
rect 17129 15991 17187 15997
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 16390 15920 16396 15972
rect 16448 15960 16454 15972
rect 17589 15963 17647 15969
rect 17589 15960 17601 15963
rect 16448 15932 17601 15960
rect 16448 15920 16454 15932
rect 17589 15929 17601 15932
rect 17635 15929 17647 15963
rect 17589 15923 17647 15929
rect 16850 15892 16856 15904
rect 12584 15864 16068 15892
rect 16811 15864 16856 15892
rect 12584 15852 12590 15864
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 1104 15802 18860 15824
rect 1104 15750 3169 15802
rect 3221 15750 3233 15802
rect 3285 15750 3297 15802
rect 3349 15750 3361 15802
rect 3413 15750 3425 15802
rect 3477 15750 7608 15802
rect 7660 15750 7672 15802
rect 7724 15750 7736 15802
rect 7788 15750 7800 15802
rect 7852 15750 7864 15802
rect 7916 15750 12047 15802
rect 12099 15750 12111 15802
rect 12163 15750 12175 15802
rect 12227 15750 12239 15802
rect 12291 15750 12303 15802
rect 12355 15750 16486 15802
rect 16538 15750 16550 15802
rect 16602 15750 16614 15802
rect 16666 15750 16678 15802
rect 16730 15750 16742 15802
rect 16794 15750 18860 15802
rect 1104 15728 18860 15750
rect 2225 15691 2283 15697
rect 2225 15657 2237 15691
rect 2271 15688 2283 15691
rect 2774 15688 2780 15700
rect 2271 15660 2780 15688
rect 2271 15657 2283 15660
rect 2225 15651 2283 15657
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 6178 15688 6184 15700
rect 6139 15660 6184 15688
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6638 15688 6644 15700
rect 6599 15660 6644 15688
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 7098 15688 7104 15700
rect 6880 15660 7104 15688
rect 6880 15648 6886 15660
rect 7098 15648 7104 15660
rect 7156 15648 7162 15700
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 8018 15688 8024 15700
rect 7248 15660 8024 15688
rect 7248 15648 7254 15660
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 9309 15691 9367 15697
rect 9309 15657 9321 15691
rect 9355 15688 9367 15691
rect 11238 15688 11244 15700
rect 9355 15660 11244 15688
rect 9355 15657 9367 15660
rect 9309 15651 9367 15657
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 15562 15688 15568 15700
rect 12492 15660 15568 15688
rect 12492 15648 12498 15660
rect 15562 15648 15568 15660
rect 15620 15648 15626 15700
rect 5166 15580 5172 15632
rect 5224 15620 5230 15632
rect 7208 15620 7236 15648
rect 5224 15592 7236 15620
rect 5224 15580 5230 15592
rect 7374 15580 7380 15632
rect 7432 15620 7438 15632
rect 7561 15623 7619 15629
rect 7561 15620 7573 15623
rect 7432 15592 7573 15620
rect 7432 15580 7438 15592
rect 7561 15589 7573 15592
rect 7607 15589 7619 15623
rect 7561 15583 7619 15589
rect 8389 15623 8447 15629
rect 8389 15589 8401 15623
rect 8435 15620 8447 15623
rect 8478 15620 8484 15632
rect 8435 15592 8484 15620
rect 8435 15589 8447 15592
rect 8389 15583 8447 15589
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 8662 15580 8668 15632
rect 8720 15620 8726 15632
rect 9766 15620 9772 15632
rect 8720 15592 9772 15620
rect 8720 15580 8726 15592
rect 9766 15580 9772 15592
rect 9824 15580 9830 15632
rect 11146 15580 11152 15632
rect 11204 15620 11210 15632
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 11204 15592 11529 15620
rect 11204 15580 11210 15592
rect 11517 15589 11529 15592
rect 11563 15589 11575 15623
rect 11517 15583 11575 15589
rect 11790 15580 11796 15632
rect 11848 15620 11854 15632
rect 11977 15623 12035 15629
rect 11977 15620 11989 15623
rect 11848 15592 11989 15620
rect 11848 15580 11854 15592
rect 11977 15589 11989 15592
rect 12023 15589 12035 15623
rect 11977 15583 12035 15589
rect 6730 15552 6736 15564
rect 6643 15524 6736 15552
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 6656 15493 6684 15524
rect 6730 15512 6736 15524
rect 6788 15552 6794 15564
rect 9214 15552 9220 15564
rect 6788 15524 9220 15552
rect 6788 15512 6794 15524
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9732 15524 10057 15552
rect 9732 15512 9738 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 10778 15512 10784 15564
rect 10836 15552 10842 15564
rect 12986 15552 12992 15564
rect 10836 15524 12992 15552
rect 10836 15512 10842 15524
rect 6641 15487 6699 15493
rect 6641 15453 6653 15487
rect 6687 15453 6699 15487
rect 6641 15447 6699 15453
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 6730 15376 6736 15428
rect 6788 15416 6794 15428
rect 6840 15416 6868 15447
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 7156 15456 7297 15484
rect 7156 15444 7162 15456
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 7285 15447 7343 15453
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15484 7619 15487
rect 8018 15484 8024 15496
rect 7607 15456 8024 15484
rect 7607 15453 7619 15456
rect 7561 15447 7619 15453
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 8159 15456 8616 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 6788 15388 6868 15416
rect 8588 15416 8616 15456
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9456 15456 9781 15484
rect 9456 15444 9462 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 11164 15470 11192 15524
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 13449 15555 13507 15561
rect 13449 15521 13461 15555
rect 13495 15552 13507 15555
rect 14550 15552 14556 15564
rect 13495 15524 14556 15552
rect 13495 15521 13507 15524
rect 13449 15515 13507 15521
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 15010 15512 15016 15564
rect 15068 15552 15074 15564
rect 18322 15552 18328 15564
rect 15068 15524 18328 15552
rect 15068 15512 15074 15524
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 13725 15487 13783 15493
rect 9769 15447 9827 15453
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 13814 15484 13820 15496
rect 13771 15456 13820 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 14323 15487 14381 15493
rect 14323 15453 14335 15487
rect 14369 15484 14381 15487
rect 14826 15484 14832 15496
rect 14369 15456 14832 15484
rect 14369 15453 14381 15456
rect 14323 15447 14381 15453
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 15746 15484 15752 15496
rect 15707 15456 15752 15484
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 16114 15484 16120 15496
rect 16075 15456 16120 15484
rect 16114 15444 16120 15456
rect 16172 15484 16178 15496
rect 16577 15487 16635 15493
rect 16577 15484 16589 15487
rect 16172 15456 16589 15484
rect 16172 15444 16178 15456
rect 16577 15453 16589 15456
rect 16623 15453 16635 15487
rect 16577 15447 16635 15453
rect 8588 15388 10272 15416
rect 13018 15388 13124 15416
rect 6788 15376 6794 15388
rect 8573 15351 8631 15357
rect 8573 15317 8585 15351
rect 8619 15348 8631 15351
rect 8846 15348 8852 15360
rect 8619 15320 8852 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 9030 15308 9036 15360
rect 9088 15348 9094 15360
rect 9674 15348 9680 15360
rect 9088 15320 9680 15348
rect 9088 15308 9094 15320
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 10244 15348 10272 15388
rect 12618 15348 12624 15360
rect 10244 15320 12624 15348
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 13096 15348 13124 15388
rect 13170 15376 13176 15428
rect 13228 15416 13234 15428
rect 13228 15388 14228 15416
rect 13228 15376 13234 15388
rect 13998 15348 14004 15360
rect 13096 15320 14004 15348
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 14200 15348 14228 15388
rect 15010 15376 15016 15428
rect 15068 15376 15074 15428
rect 16853 15419 16911 15425
rect 16853 15385 16865 15419
rect 16899 15385 16911 15419
rect 16853 15379 16911 15385
rect 16868 15348 16896 15379
rect 17310 15376 17316 15428
rect 17368 15376 17374 15428
rect 14200 15320 16896 15348
rect 18325 15351 18383 15357
rect 18325 15317 18337 15351
rect 18371 15348 18383 15351
rect 18414 15348 18420 15360
rect 18371 15320 18420 15348
rect 18371 15317 18383 15320
rect 18325 15311 18383 15317
rect 18414 15308 18420 15320
rect 18472 15308 18478 15360
rect 1104 15258 19019 15280
rect 1104 15206 5388 15258
rect 5440 15206 5452 15258
rect 5504 15206 5516 15258
rect 5568 15206 5580 15258
rect 5632 15206 5644 15258
rect 5696 15206 9827 15258
rect 9879 15206 9891 15258
rect 9943 15206 9955 15258
rect 10007 15206 10019 15258
rect 10071 15206 10083 15258
rect 10135 15206 14266 15258
rect 14318 15206 14330 15258
rect 14382 15206 14394 15258
rect 14446 15206 14458 15258
rect 14510 15206 14522 15258
rect 14574 15206 18705 15258
rect 18757 15206 18769 15258
rect 18821 15206 18833 15258
rect 18885 15206 18897 15258
rect 18949 15206 18961 15258
rect 19013 15206 19019 15258
rect 1104 15184 19019 15206
rect 7926 15144 7932 15156
rect 7887 15116 7932 15144
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 9033 15147 9091 15153
rect 9033 15113 9045 15147
rect 9079 15144 9091 15147
rect 11606 15144 11612 15156
rect 9079 15116 11612 15144
rect 9079 15113 9091 15116
rect 9033 15107 9091 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 12526 15144 12532 15156
rect 12487 15116 12532 15144
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12894 15144 12900 15156
rect 12676 15116 12900 15144
rect 12676 15104 12682 15116
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 12989 15147 13047 15153
rect 12989 15113 13001 15147
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 8665 15079 8723 15085
rect 8665 15045 8677 15079
rect 8711 15076 8723 15079
rect 12434 15076 12440 15088
rect 8711 15048 10732 15076
rect 8711 15045 8723 15048
rect 8665 15039 8723 15045
rect 1486 14968 1492 15020
rect 1544 15008 1550 15020
rect 1581 15011 1639 15017
rect 1581 15008 1593 15011
rect 1544 14980 1593 15008
rect 1544 14968 1550 14980
rect 1581 14977 1593 14980
rect 1627 14977 1639 15011
rect 7190 15008 7196 15020
rect 7151 14980 7196 15008
rect 1581 14971 1639 14977
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 8110 15008 8116 15020
rect 8071 14980 8116 15008
rect 7377 14971 7435 14977
rect 7392 14940 7420 14971
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 8573 15011 8631 15017
rect 8573 14977 8585 15011
rect 8619 14977 8631 15011
rect 8846 15008 8852 15020
rect 8807 14980 8852 15008
rect 8573 14971 8631 14977
rect 7300 14912 7420 14940
rect 6733 14807 6791 14813
rect 6733 14773 6745 14807
rect 6779 14804 6791 14807
rect 6822 14804 6828 14816
rect 6779 14776 6828 14804
rect 6779 14773 6791 14776
rect 6733 14767 6791 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7300 14804 7328 14912
rect 7377 14875 7435 14881
rect 7377 14841 7389 14875
rect 7423 14872 7435 14875
rect 8588 14872 8616 14971
rect 8846 14968 8852 14980
rect 8904 14968 8910 15020
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 15008 9735 15011
rect 10410 15008 10416 15020
rect 9723 14980 10416 15008
rect 9723 14977 9735 14980
rect 9677 14971 9735 14977
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 10594 15008 10600 15020
rect 10551 14980 10600 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 9640 14912 9781 14940
rect 9640 14900 9646 14912
rect 9769 14909 9781 14912
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14940 10103 14943
rect 10318 14940 10324 14952
rect 10091 14912 10324 14940
rect 10091 14909 10103 14912
rect 10045 14903 10103 14909
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 10226 14872 10232 14884
rect 7423 14844 10232 14872
rect 7423 14841 7435 14844
rect 7377 14835 7435 14841
rect 10226 14832 10232 14844
rect 10284 14832 10290 14884
rect 10704 14872 10732 15048
rect 10888 15048 12440 15076
rect 10778 14968 10784 15020
rect 10836 15008 10842 15020
rect 10888 15017 10916 15048
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 13004 15076 13032 15107
rect 13538 15104 13544 15156
rect 13596 15144 13602 15156
rect 13814 15144 13820 15156
rect 13596 15116 13820 15144
rect 13596 15104 13602 15116
rect 13814 15104 13820 15116
rect 13872 15144 13878 15156
rect 13872 15116 15056 15144
rect 13872 15104 13878 15116
rect 14366 15076 14372 15088
rect 12728 15048 13032 15076
rect 14030 15048 14372 15076
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 10836 14980 10885 15008
rect 10836 14968 10842 14980
rect 10873 14977 10885 14980
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 11112 14980 12173 15008
rect 11112 14968 11118 14980
rect 12161 14977 12173 14980
rect 12207 15008 12219 15011
rect 12728 15008 12756 15048
rect 14366 15036 14372 15048
rect 14424 15036 14430 15088
rect 14461 15079 14519 15085
rect 14461 15045 14473 15079
rect 14507 15076 14519 15079
rect 14918 15076 14924 15088
rect 14507 15048 14924 15076
rect 14507 15045 14519 15048
rect 14461 15039 14519 15045
rect 14918 15036 14924 15048
rect 14976 15036 14982 15088
rect 15028 15020 15056 15116
rect 15470 15104 15476 15156
rect 15528 15144 15534 15156
rect 17862 15144 17868 15156
rect 15528 15116 17868 15144
rect 15528 15104 15534 15116
rect 17862 15104 17868 15116
rect 17920 15144 17926 15156
rect 17920 15116 18092 15144
rect 17920 15104 17926 15116
rect 15933 15079 15991 15085
rect 15933 15045 15945 15079
rect 15979 15076 15991 15079
rect 17218 15076 17224 15088
rect 15979 15048 17224 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 17218 15036 17224 15048
rect 17276 15076 17282 15088
rect 17954 15076 17960 15088
rect 17276 15048 17960 15076
rect 17276 15036 17282 15048
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 18064 15085 18092 15116
rect 18049 15079 18107 15085
rect 18049 15045 18061 15079
rect 18095 15045 18107 15079
rect 18049 15039 18107 15045
rect 12207 14980 12756 15008
rect 14737 15011 14795 15017
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 14737 14977 14749 15011
rect 14783 15008 14795 15011
rect 15010 15008 15016 15020
rect 14783 14980 15016 15008
rect 14783 14977 14795 14980
rect 14737 14971 14795 14977
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 17405 15011 17463 15017
rect 17405 14977 17417 15011
rect 17451 15008 17463 15011
rect 17770 15008 17776 15020
rect 17451 14980 17776 15008
rect 17451 14977 17463 14980
rect 17405 14971 17463 14977
rect 17770 14968 17776 14980
rect 17828 14968 17834 15020
rect 18230 15008 18236 15020
rect 18191 14980 18236 15008
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18380 14980 18425 15008
rect 18380 14968 18386 14980
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14940 11023 14943
rect 11698 14940 11704 14952
rect 11011 14912 11704 14940
rect 11011 14909 11023 14912
rect 10965 14903 11023 14909
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 11882 14940 11888 14952
rect 11843 14912 11888 14940
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 12069 14943 12127 14949
rect 12069 14909 12081 14943
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 10704 14844 11284 14872
rect 9030 14804 9036 14816
rect 7300 14776 9036 14804
rect 9030 14764 9036 14776
rect 9088 14764 9094 14816
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 10778 14804 10784 14816
rect 10100 14776 10784 14804
rect 10100 14764 10106 14776
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11146 14804 11152 14816
rect 11107 14776 11152 14804
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11256 14804 11284 14844
rect 11514 14832 11520 14884
rect 11572 14872 11578 14884
rect 12084 14872 12112 14903
rect 12986 14900 12992 14952
rect 13044 14940 13050 14952
rect 15381 14943 15439 14949
rect 13044 14912 14688 14940
rect 13044 14900 13050 14912
rect 11572 14844 12112 14872
rect 14660 14872 14688 14912
rect 15381 14909 15393 14943
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 15473 14943 15531 14949
rect 15473 14909 15485 14943
rect 15519 14940 15531 14943
rect 16114 14940 16120 14952
rect 15519 14912 16120 14940
rect 15519 14909 15531 14912
rect 15473 14903 15531 14909
rect 15286 14872 15292 14884
rect 14660 14844 15292 14872
rect 11572 14832 11578 14844
rect 15286 14832 15292 14844
rect 15344 14832 15350 14884
rect 13078 14804 13084 14816
rect 11256 14776 13084 14804
rect 13078 14764 13084 14776
rect 13136 14804 13142 14816
rect 15197 14807 15255 14813
rect 15197 14804 15209 14807
rect 13136 14776 15209 14804
rect 13136 14764 13142 14776
rect 15197 14773 15209 14776
rect 15243 14773 15255 14807
rect 15396 14804 15424 14903
rect 16114 14900 16120 14912
rect 16172 14940 16178 14952
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 16172 14912 16865 14940
rect 16172 14900 16178 14912
rect 16853 14909 16865 14912
rect 16899 14940 16911 14943
rect 17034 14940 17040 14952
rect 16899 14912 17040 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 17126 14900 17132 14952
rect 17184 14940 17190 14952
rect 17494 14940 17500 14952
rect 17184 14912 17229 14940
rect 17455 14912 17500 14940
rect 17184 14900 17190 14912
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 15933 14875 15991 14881
rect 15933 14841 15945 14875
rect 15979 14872 15991 14875
rect 16390 14872 16396 14884
rect 15979 14844 16396 14872
rect 15979 14841 15991 14844
rect 15933 14835 15991 14841
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 17678 14804 17684 14816
rect 15396 14776 17684 14804
rect 15197 14767 15255 14773
rect 17678 14764 17684 14776
rect 17736 14764 17742 14816
rect 18046 14804 18052 14816
rect 18007 14776 18052 14804
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 1104 14714 18860 14736
rect 1104 14662 3169 14714
rect 3221 14662 3233 14714
rect 3285 14662 3297 14714
rect 3349 14662 3361 14714
rect 3413 14662 3425 14714
rect 3477 14662 7608 14714
rect 7660 14662 7672 14714
rect 7724 14662 7736 14714
rect 7788 14662 7800 14714
rect 7852 14662 7864 14714
rect 7916 14662 12047 14714
rect 12099 14662 12111 14714
rect 12163 14662 12175 14714
rect 12227 14662 12239 14714
rect 12291 14662 12303 14714
rect 12355 14662 16486 14714
rect 16538 14662 16550 14714
rect 16602 14662 16614 14714
rect 16666 14662 16678 14714
rect 16730 14662 16742 14714
rect 16794 14662 18860 14714
rect 1104 14640 18860 14662
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 7101 14603 7159 14609
rect 7101 14600 7113 14603
rect 7064 14572 7113 14600
rect 7064 14560 7070 14572
rect 7101 14569 7113 14572
rect 7147 14569 7159 14603
rect 7926 14600 7932 14612
rect 7887 14572 7932 14600
rect 7101 14563 7159 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8570 14600 8576 14612
rect 8531 14572 8576 14600
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 9401 14603 9459 14609
rect 9401 14569 9413 14603
rect 9447 14600 9459 14603
rect 10318 14600 10324 14612
rect 9447 14572 10324 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 11514 14600 11520 14612
rect 11475 14572 11520 14600
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 11698 14560 11704 14612
rect 11756 14600 11762 14612
rect 15654 14600 15660 14612
rect 11756 14572 15660 14600
rect 11756 14560 11762 14572
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 8202 14492 8208 14544
rect 8260 14532 8266 14544
rect 10134 14532 10140 14544
rect 8260 14504 10140 14532
rect 8260 14492 8266 14504
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 10505 14535 10563 14541
rect 10505 14501 10517 14535
rect 10551 14532 10563 14535
rect 11422 14532 11428 14544
rect 10551 14504 11428 14532
rect 10551 14501 10563 14504
rect 10505 14495 10563 14501
rect 11422 14492 11428 14504
rect 11480 14492 11486 14544
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10594 14464 10600 14476
rect 10091 14436 10600 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 11241 14467 11299 14473
rect 11241 14433 11253 14467
rect 11287 14464 11299 14467
rect 11514 14464 11520 14476
rect 11287 14436 11520 14464
rect 11287 14433 11299 14436
rect 11241 14427 11299 14433
rect 11514 14424 11520 14436
rect 11572 14464 11578 14476
rect 11790 14464 11796 14476
rect 11572 14436 11796 14464
rect 11572 14424 11578 14436
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 13446 14464 13452 14476
rect 11900 14436 13452 14464
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 8386 14396 8392 14408
rect 8347 14368 8392 14396
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 10321 14399 10379 14405
rect 9232 14368 10272 14396
rect 7190 14288 7196 14340
rect 7248 14328 7254 14340
rect 9232 14337 9260 14368
rect 9217 14331 9275 14337
rect 9217 14328 9229 14331
rect 7248 14300 9229 14328
rect 7248 14288 7254 14300
rect 9217 14297 9229 14300
rect 9263 14297 9275 14331
rect 9217 14291 9275 14297
rect 9433 14331 9491 14337
rect 9433 14297 9445 14331
rect 9479 14328 9491 14331
rect 10042 14328 10048 14340
rect 9479 14300 10048 14328
rect 9479 14297 9491 14300
rect 9433 14291 9491 14297
rect 10042 14288 10048 14300
rect 10100 14288 10106 14340
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 9582 14260 9588 14272
rect 8352 14232 9588 14260
rect 8352 14220 8358 14232
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 10244 14260 10272 14368
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10778 14396 10784 14408
rect 10367 14368 10784 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 11112 14368 11161 14396
rect 11112 14356 11118 14368
rect 11149 14365 11161 14368
rect 11195 14396 11207 14399
rect 11900 14396 11928 14436
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 13725 14467 13783 14473
rect 13725 14433 13737 14467
rect 13771 14464 13783 14467
rect 13906 14464 13912 14476
rect 13771 14436 13912 14464
rect 13771 14433 13783 14436
rect 13725 14427 13783 14433
rect 13906 14424 13912 14436
rect 13964 14464 13970 14476
rect 14277 14467 14335 14473
rect 14277 14464 14289 14467
rect 13964 14436 14289 14464
rect 13964 14424 13970 14436
rect 14277 14433 14289 14436
rect 14323 14433 14335 14467
rect 14277 14427 14335 14433
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 14642 14464 14648 14476
rect 14599 14436 14648 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 16485 14467 16543 14473
rect 16485 14464 16497 14467
rect 15068 14436 16497 14464
rect 15068 14424 15074 14436
rect 16485 14433 16497 14436
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 17402 14424 17408 14476
rect 17460 14464 17466 14476
rect 17770 14464 17776 14476
rect 17460 14436 17776 14464
rect 17460 14424 17466 14436
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 18012 14436 18245 14464
rect 18012 14424 18018 14436
rect 18233 14433 18245 14436
rect 18279 14433 18291 14467
rect 18233 14427 18291 14433
rect 11195 14368 11928 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11238 14288 11244 14340
rect 11296 14328 11302 14340
rect 11422 14328 11428 14340
rect 11296 14300 11428 14328
rect 11296 14288 11302 14300
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 12986 14288 12992 14340
rect 13044 14288 13050 14340
rect 13449 14331 13507 14337
rect 13449 14297 13461 14331
rect 13495 14328 13507 14331
rect 13906 14328 13912 14340
rect 13495 14300 13912 14328
rect 13495 14297 13507 14300
rect 13449 14291 13507 14297
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 15286 14288 15292 14340
rect 15344 14288 15350 14340
rect 16206 14328 16212 14340
rect 15948 14300 16212 14328
rect 11698 14260 11704 14272
rect 10244 14232 11704 14260
rect 11698 14220 11704 14232
rect 11756 14260 11762 14272
rect 11974 14260 11980 14272
rect 11756 14232 11980 14260
rect 11756 14220 11762 14232
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 15948 14260 15976 14300
rect 16206 14288 16212 14300
rect 16264 14288 16270 14340
rect 16761 14331 16819 14337
rect 16761 14297 16773 14331
rect 16807 14328 16819 14331
rect 16850 14328 16856 14340
rect 16807 14300 16856 14328
rect 16807 14297 16819 14300
rect 16761 14291 16819 14297
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 17770 14288 17776 14340
rect 17828 14288 17834 14340
rect 13136 14232 15976 14260
rect 16025 14263 16083 14269
rect 13136 14220 13142 14232
rect 16025 14229 16037 14263
rect 16071 14260 16083 14263
rect 17678 14260 17684 14272
rect 16071 14232 17684 14260
rect 16071 14229 16083 14232
rect 16025 14223 16083 14229
rect 17678 14220 17684 14232
rect 17736 14220 17742 14272
rect 1104 14170 19019 14192
rect 1104 14118 5388 14170
rect 5440 14118 5452 14170
rect 5504 14118 5516 14170
rect 5568 14118 5580 14170
rect 5632 14118 5644 14170
rect 5696 14118 9827 14170
rect 9879 14118 9891 14170
rect 9943 14118 9955 14170
rect 10007 14118 10019 14170
rect 10071 14118 10083 14170
rect 10135 14118 14266 14170
rect 14318 14118 14330 14170
rect 14382 14118 14394 14170
rect 14446 14118 14458 14170
rect 14510 14118 14522 14170
rect 14574 14118 18705 14170
rect 18757 14118 18769 14170
rect 18821 14118 18833 14170
rect 18885 14118 18897 14170
rect 18949 14118 18961 14170
rect 19013 14118 19019 14170
rect 1104 14096 19019 14118
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 12618 14056 12624 14068
rect 9640 14028 12624 14056
rect 9640 14016 9646 14028
rect 9309 13991 9367 13997
rect 9309 13957 9321 13991
rect 9355 13988 9367 13991
rect 10502 13988 10508 14000
rect 9355 13960 10508 13988
rect 9355 13957 9367 13960
rect 9309 13951 9367 13957
rect 10502 13948 10508 13960
rect 10560 13948 10566 14000
rect 10965 13991 11023 13997
rect 10965 13957 10977 13991
rect 11011 13988 11023 13991
rect 11238 13988 11244 14000
rect 11011 13960 11244 13988
rect 11011 13957 11023 13960
rect 10965 13951 11023 13957
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 8754 13920 8760 13932
rect 8715 13892 8760 13920
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9398 13920 9404 13932
rect 9359 13892 9404 13920
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10042 13920 10048 13932
rect 9732 13892 10048 13920
rect 9732 13880 9738 13892
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10594 13880 10600 13932
rect 10652 13920 10658 13932
rect 10689 13923 10747 13929
rect 10689 13920 10701 13923
rect 10652 13892 10701 13920
rect 10652 13880 10658 13892
rect 10689 13889 10701 13892
rect 10735 13889 10747 13923
rect 10870 13920 10876 13932
rect 10831 13892 10876 13920
rect 10689 13883 10747 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 11062 13923 11120 13929
rect 11062 13889 11074 13923
rect 11108 13920 11120 13923
rect 11348 13920 11376 14028
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 12894 14056 12900 14068
rect 12807 14028 12900 14056
rect 12894 14016 12900 14028
rect 12952 14056 12958 14068
rect 13078 14056 13084 14068
rect 12952 14028 13084 14056
rect 12952 14016 12958 14028
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13280 14028 15056 14056
rect 11974 13948 11980 14000
rect 12032 13988 12038 14000
rect 12738 13991 12796 13997
rect 12738 13988 12750 13991
rect 12032 13960 12750 13988
rect 12032 13948 12038 13960
rect 12738 13957 12750 13960
rect 12784 13988 12796 13991
rect 12986 13988 12992 14000
rect 12784 13960 12992 13988
rect 12784 13957 12796 13960
rect 12738 13951 12796 13957
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 12250 13929 12256 13932
rect 11108 13892 11376 13920
rect 12241 13923 12256 13929
rect 11108 13889 11120 13892
rect 11062 13883 11120 13889
rect 12241 13889 12253 13923
rect 12241 13883 12256 13889
rect 12250 13880 12256 13883
rect 12308 13880 12314 13932
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 12894 13920 12900 13932
rect 12667 13892 12900 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 7340 13824 9873 13852
rect 7340 13812 7346 13824
rect 9861 13821 9873 13824
rect 9907 13852 9919 13855
rect 10318 13852 10324 13864
rect 9907 13824 10324 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 11238 13812 11244 13864
rect 11296 13852 11302 13864
rect 12529 13855 12587 13861
rect 12529 13852 12541 13855
rect 11296 13824 12541 13852
rect 11296 13812 11302 13824
rect 12529 13821 12541 13824
rect 12575 13852 12587 13855
rect 13280 13852 13308 14028
rect 13538 13988 13544 14000
rect 13372 13960 13544 13988
rect 13372 13929 13400 13960
rect 13538 13948 13544 13960
rect 13596 13948 13602 14000
rect 14918 13988 14924 14000
rect 14858 13960 14924 13988
rect 14918 13948 14924 13960
rect 14976 13948 14982 14000
rect 15028 13988 15056 14028
rect 15102 14016 15108 14068
rect 15160 14056 15166 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 15160 14028 16865 14056
rect 15160 14016 15166 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 18115 14059 18173 14065
rect 18115 14056 18127 14059
rect 16853 14019 16911 14025
rect 16960 14028 18127 14056
rect 15194 13988 15200 14000
rect 15028 13960 15200 13988
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 15933 13991 15991 13997
rect 15933 13988 15945 13991
rect 15304 13960 15945 13988
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 15304 13920 15332 13960
rect 15933 13957 15945 13960
rect 15979 13957 15991 13991
rect 15933 13951 15991 13957
rect 16022 13948 16028 14000
rect 16080 13997 16086 14000
rect 16080 13991 16109 13997
rect 16097 13957 16109 13991
rect 16960 13988 16988 14028
rect 18115 14025 18127 14028
rect 18161 14025 18173 14059
rect 18115 14019 18173 14025
rect 16080 13951 16109 13957
rect 16500 13960 16988 13988
rect 16080 13948 16086 13951
rect 13357 13883 13415 13889
rect 14844 13892 15332 13920
rect 13633 13855 13691 13861
rect 13633 13852 13645 13855
rect 12575 13824 13308 13852
rect 13372 13824 13645 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 7466 13744 7472 13796
rect 7524 13784 7530 13796
rect 13372 13784 13400 13824
rect 13633 13821 13645 13824
rect 13679 13821 13691 13855
rect 13633 13815 13691 13821
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14642 13852 14648 13864
rect 14056 13824 14648 13852
rect 14056 13812 14062 13824
rect 14642 13812 14648 13824
rect 14700 13852 14706 13864
rect 14844 13852 14872 13892
rect 15562 13880 15568 13932
rect 15620 13920 15626 13932
rect 15749 13923 15807 13929
rect 15620 13892 15665 13920
rect 15620 13880 15626 13892
rect 15749 13889 15761 13923
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 14700 13824 14872 13852
rect 14700 13812 14706 13824
rect 15654 13812 15660 13864
rect 15712 13852 15718 13864
rect 15764 13852 15792 13883
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 15896 13892 15941 13920
rect 15896 13880 15902 13892
rect 15712 13824 15792 13852
rect 15712 13812 15718 13824
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 16264 13824 16309 13852
rect 16264 13812 16270 13824
rect 15378 13784 15384 13796
rect 7524 13756 13400 13784
rect 15120 13756 15384 13784
rect 7524 13744 7530 13756
rect 15120 13728 15148 13756
rect 15378 13744 15384 13756
rect 15436 13784 15442 13796
rect 16500 13784 16528 13960
rect 17862 13948 17868 14000
rect 17920 13988 17926 14000
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 17920 13960 18337 13988
rect 17920 13948 17926 13960
rect 18325 13957 18337 13960
rect 18371 13957 18383 13991
rect 18325 13951 18383 13957
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17218 13920 17224 13932
rect 17083 13892 17224 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 17310 13880 17316 13932
rect 17368 13920 17374 13932
rect 17497 13923 17555 13929
rect 17497 13920 17509 13923
rect 17368 13892 17509 13920
rect 17368 13880 17374 13892
rect 17497 13889 17509 13892
rect 17543 13889 17555 13923
rect 17497 13883 17555 13889
rect 17126 13852 17132 13864
rect 17087 13824 17132 13852
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 18414 13784 18420 13796
rect 15436 13756 16528 13784
rect 17420 13756 18420 13784
rect 15436 13744 15442 13756
rect 10229 13719 10287 13725
rect 10229 13685 10241 13719
rect 10275 13716 10287 13719
rect 10318 13716 10324 13728
rect 10275 13688 10324 13716
rect 10275 13685 10287 13688
rect 10229 13679 10287 13685
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 10689 13719 10747 13725
rect 10689 13716 10701 13719
rect 10560 13688 10701 13716
rect 10560 13676 10566 13688
rect 10689 13685 10701 13688
rect 10735 13685 10747 13719
rect 10689 13679 10747 13685
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 11790 13716 11796 13728
rect 11296 13688 11796 13716
rect 11296 13676 11302 13688
rect 11790 13676 11796 13688
rect 11848 13716 11854 13728
rect 13354 13716 13360 13728
rect 11848 13688 13360 13716
rect 11848 13676 11854 13688
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 15102 13716 15108 13728
rect 15063 13688 15108 13716
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 17034 13676 17040 13728
rect 17092 13716 17098 13728
rect 17420 13725 17448 13756
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 17405 13719 17463 13725
rect 17405 13716 17417 13719
rect 17092 13688 17417 13716
rect 17092 13676 17098 13688
rect 17405 13685 17417 13688
rect 17451 13685 17463 13719
rect 17954 13716 17960 13728
rect 17915 13688 17960 13716
rect 17405 13679 17463 13685
rect 17954 13676 17960 13688
rect 18012 13676 18018 13728
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 18141 13719 18199 13725
rect 18141 13716 18153 13719
rect 18104 13688 18153 13716
rect 18104 13676 18110 13688
rect 18141 13685 18153 13688
rect 18187 13716 18199 13719
rect 18230 13716 18236 13728
rect 18187 13688 18236 13716
rect 18187 13685 18199 13688
rect 18141 13679 18199 13685
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 1104 13626 18860 13648
rect 1104 13574 3169 13626
rect 3221 13574 3233 13626
rect 3285 13574 3297 13626
rect 3349 13574 3361 13626
rect 3413 13574 3425 13626
rect 3477 13574 7608 13626
rect 7660 13574 7672 13626
rect 7724 13574 7736 13626
rect 7788 13574 7800 13626
rect 7852 13574 7864 13626
rect 7916 13574 12047 13626
rect 12099 13574 12111 13626
rect 12163 13574 12175 13626
rect 12227 13574 12239 13626
rect 12291 13574 12303 13626
rect 12355 13574 16486 13626
rect 16538 13574 16550 13626
rect 16602 13574 16614 13626
rect 16666 13574 16678 13626
rect 16730 13574 16742 13626
rect 16794 13574 18860 13626
rect 1104 13552 18860 13574
rect 9953 13515 10011 13521
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 11054 13512 11060 13524
rect 9999 13484 11060 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 11164 13484 12112 13512
rect 10502 13444 10508 13456
rect 10428 13416 10508 13444
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 10428 13376 10456 13416
rect 10502 13404 10508 13416
rect 10560 13404 10566 13456
rect 10597 13447 10655 13453
rect 10597 13413 10609 13447
rect 10643 13444 10655 13447
rect 11164 13444 11192 13484
rect 10643 13416 11192 13444
rect 10643 13413 10655 13416
rect 10597 13407 10655 13413
rect 11238 13404 11244 13456
rect 11296 13404 11302 13456
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 11974 13444 11980 13456
rect 11664 13416 11980 13444
rect 11664 13404 11670 13416
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 12084 13444 12112 13484
rect 12158 13472 12164 13524
rect 12216 13512 12222 13524
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 12216 13484 12265 13512
rect 12216 13472 12222 13484
rect 12253 13481 12265 13484
rect 12299 13481 12311 13515
rect 16022 13512 16028 13524
rect 12253 13475 12311 13481
rect 12452 13484 16028 13512
rect 12452 13444 12480 13484
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 17034 13512 17040 13524
rect 16995 13484 17040 13512
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 17589 13515 17647 13521
rect 17589 13512 17601 13515
rect 17552 13484 17601 13512
rect 17552 13472 17558 13484
rect 17589 13481 17601 13484
rect 17635 13481 17647 13515
rect 17862 13512 17868 13524
rect 17823 13484 17868 13512
rect 17589 13475 17647 13481
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 12084 13416 12480 13444
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 13722 13444 13728 13456
rect 12584 13416 13728 13444
rect 12584 13404 12590 13416
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 16408 13416 17908 13444
rect 11256 13376 11284 13404
rect 16408 13388 16436 13416
rect 17512 13388 17540 13416
rect 6788 13348 10456 13376
rect 6788 13336 6794 13348
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 7098 13268 7104 13320
rect 7156 13308 7162 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 7156 13280 9781 13308
rect 7156 13268 7162 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 9784 13240 9812 13271
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 10428 13317 10456 13348
rect 10704 13348 11284 13376
rect 11333 13379 11391 13385
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 9916 13280 9965 13308
rect 9916 13268 9922 13280
rect 9953 13277 9965 13280
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 10594 13308 10600 13320
rect 10551 13280 10600 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 10704 13317 10732 13348
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 13081 13379 13139 13385
rect 11379 13348 13032 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 11146 13308 11152 13320
rect 11107 13280 11152 13308
rect 10689 13271 10747 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 11238 13268 11244 13320
rect 11296 13310 11302 13320
rect 11471 13311 11529 13317
rect 11296 13308 11376 13310
rect 11471 13308 11483 13311
rect 11296 13282 11483 13308
rect 11296 13268 11302 13282
rect 11348 13280 11483 13282
rect 11471 13277 11483 13280
rect 11517 13277 11529 13311
rect 11471 13271 11529 13277
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 11664 13280 11709 13308
rect 11664 13268 11670 13280
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 11992 13308 12296 13310
rect 12618 13308 12624 13320
rect 11940 13282 12296 13308
rect 11940 13280 12020 13282
rect 11940 13268 11946 13280
rect 11624 13240 11652 13268
rect 12268 13249 12296 13282
rect 12579 13280 12624 13308
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 13004 13308 13032 13348
rect 13081 13345 13093 13379
rect 13127 13376 13139 13379
rect 13170 13376 13176 13388
rect 13127 13348 13176 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 13354 13376 13360 13388
rect 13315 13348 13360 13376
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 13446 13336 13452 13388
rect 13504 13376 13510 13388
rect 16298 13376 16304 13388
rect 13504 13348 16304 13376
rect 13504 13336 13510 13348
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 16390 13336 16396 13388
rect 16448 13336 16454 13388
rect 17310 13376 17316 13388
rect 16776 13348 17316 13376
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 13004 13280 13277 13308
rect 13265 13277 13277 13280
rect 13311 13308 13323 13311
rect 13538 13308 13544 13320
rect 13311 13280 13544 13308
rect 13311 13277 13323 13280
rect 13265 13271 13323 13277
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13872 13280 14289 13308
rect 13872 13268 13878 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16408 13308 16436 13336
rect 16776 13320 16804 13348
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 17494 13336 17500 13388
rect 17552 13336 17558 13388
rect 17880 13385 17908 13416
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13345 17923 13379
rect 17865 13339 17923 13345
rect 16666 13308 16672 13320
rect 15896 13280 16436 13308
rect 16627 13280 16672 13308
rect 15896 13268 15902 13280
rect 9784 13212 11652 13240
rect 12253 13243 12311 13249
rect 12253 13209 12265 13243
rect 12299 13209 12311 13243
rect 12253 13203 12311 13209
rect 12342 13200 12348 13252
rect 12400 13240 12406 13252
rect 14553 13243 14611 13249
rect 14553 13240 14565 13243
rect 12400 13212 14565 13240
rect 12400 13200 12406 13212
rect 14553 13209 14565 13212
rect 14599 13209 14611 13243
rect 14553 13203 14611 13209
rect 15286 13200 15292 13252
rect 15344 13200 15350 13252
rect 16206 13240 16212 13252
rect 15948 13212 16212 13240
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 10410 13172 10416 13184
rect 8444 13144 10416 13172
rect 8444 13132 8450 13144
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 11241 13175 11299 13181
rect 11241 13141 11253 13175
rect 11287 13172 11299 13175
rect 11882 13172 11888 13184
rect 11287 13144 11888 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12069 13175 12127 13181
rect 12069 13172 12081 13175
rect 12032 13144 12081 13172
rect 12032 13132 12038 13144
rect 12069 13141 12081 13144
rect 12115 13141 12127 13175
rect 12069 13135 12127 13141
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12894 13172 12900 13184
rect 12492 13144 12900 13172
rect 12492 13132 12498 13144
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 13725 13175 13783 13181
rect 13725 13141 13737 13175
rect 13771 13172 13783 13175
rect 15948 13172 15976 13212
rect 16206 13200 16212 13212
rect 16264 13200 16270 13252
rect 13771 13144 15976 13172
rect 16025 13175 16083 13181
rect 13771 13141 13783 13144
rect 13725 13135 13783 13141
rect 16025 13141 16037 13175
rect 16071 13172 16083 13175
rect 16316 13172 16344 13280
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 18141 13311 18199 13317
rect 16816 13280 16861 13308
rect 16816 13268 16822 13280
rect 18141 13277 18153 13311
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 17126 13240 17132 13252
rect 16448 13212 17132 13240
rect 16448 13200 16454 13212
rect 17126 13200 17132 13212
rect 17184 13200 17190 13252
rect 17678 13200 17684 13252
rect 17736 13240 17742 13252
rect 18156 13240 18184 13271
rect 17736 13212 18184 13240
rect 17736 13200 17742 13212
rect 16482 13172 16488 13184
rect 16071 13144 16344 13172
rect 16443 13144 16488 13172
rect 16071 13141 16083 13144
rect 16025 13135 16083 13141
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 17034 13132 17040 13184
rect 17092 13172 17098 13184
rect 17862 13172 17868 13184
rect 17092 13144 17868 13172
rect 17092 13132 17098 13144
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 1104 13082 19019 13104
rect 1104 13030 5388 13082
rect 5440 13030 5452 13082
rect 5504 13030 5516 13082
rect 5568 13030 5580 13082
rect 5632 13030 5644 13082
rect 5696 13030 9827 13082
rect 9879 13030 9891 13082
rect 9943 13030 9955 13082
rect 10007 13030 10019 13082
rect 10071 13030 10083 13082
rect 10135 13030 14266 13082
rect 14318 13030 14330 13082
rect 14382 13030 14394 13082
rect 14446 13030 14458 13082
rect 14510 13030 14522 13082
rect 14574 13030 18705 13082
rect 18757 13030 18769 13082
rect 18821 13030 18833 13082
rect 18885 13030 18897 13082
rect 18949 13030 18961 13082
rect 19013 13030 19019 13082
rect 1104 13008 19019 13030
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 11146 12968 11152 12980
rect 9364 12940 11152 12968
rect 9364 12928 9370 12940
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12710 12968 12716 12980
rect 12299 12940 12716 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 14182 12968 14188 12980
rect 13320 12940 14188 12968
rect 13320 12928 13326 12940
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14918 12928 14924 12980
rect 14976 12968 14982 12980
rect 17402 12968 17408 12980
rect 14976 12940 16436 12968
rect 17363 12940 17408 12968
rect 14976 12928 14982 12940
rect 5994 12860 6000 12912
rect 6052 12900 6058 12912
rect 6052 12872 11008 12900
rect 6052 12860 6058 12872
rect 10502 12832 10508 12844
rect 10463 12804 10508 12832
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 10980 12841 11008 12872
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 14001 12903 14059 12909
rect 14001 12900 14013 12903
rect 11940 12872 14013 12900
rect 11940 12860 11946 12872
rect 14001 12869 14013 12872
rect 14047 12869 14059 12903
rect 14001 12863 14059 12869
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 16085 12903 16143 12909
rect 16085 12900 16097 12903
rect 15344 12872 16097 12900
rect 15344 12860 15350 12872
rect 16085 12869 16097 12872
rect 16131 12869 16143 12903
rect 16298 12900 16304 12912
rect 16259 12872 16304 12900
rect 16085 12863 16143 12869
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 16408 12900 16436 12940
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 16408 12872 17908 12900
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12832 11023 12835
rect 11054 12832 11060 12844
rect 11011 12804 11060 12832
rect 11011 12801 11023 12804
rect 10965 12795 11023 12801
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 9030 12656 9036 12708
rect 9088 12696 9094 12708
rect 10962 12696 10968 12708
rect 9088 12668 10640 12696
rect 10923 12668 10968 12696
rect 9088 12656 9094 12668
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 10502 12628 10508 12640
rect 8536 12600 10508 12628
rect 8536 12588 8542 12600
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 10612 12628 10640 12668
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 11164 12696 11192 12795
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11756 12804 11805 12832
rect 11756 12792 11762 12804
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 12434 12832 12440 12844
rect 12115 12804 12440 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 12526 12792 12532 12844
rect 12584 12832 12590 12844
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12584 12804 12909 12832
rect 12584 12792 12590 12804
rect 12897 12801 12909 12804
rect 12943 12832 12955 12835
rect 13078 12832 13084 12844
rect 12943 12804 13084 12832
rect 12943 12801 12955 12804
rect 12897 12795 12955 12801
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 15378 12832 15384 12844
rect 15134 12804 15384 12832
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 16390 12832 16396 12844
rect 15620 12804 16396 12832
rect 15620 12792 15626 12804
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16504 12804 16865 12832
rect 12802 12764 12808 12776
rect 12763 12736 12808 12764
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 13262 12764 13268 12776
rect 13223 12736 13268 12764
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13722 12764 13728 12776
rect 13683 12736 13728 12764
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 13832 12736 15700 12764
rect 11514 12696 11520 12708
rect 11164 12668 11520 12696
rect 11514 12656 11520 12668
rect 11572 12696 11578 12708
rect 12618 12696 12624 12708
rect 11572 12668 12624 12696
rect 11572 12656 11578 12668
rect 12618 12656 12624 12668
rect 12676 12696 12682 12708
rect 13832 12696 13860 12736
rect 12676 12668 13860 12696
rect 12676 12656 12682 12668
rect 15286 12656 15292 12708
rect 15344 12656 15350 12708
rect 11882 12628 11888 12640
rect 10612 12600 11888 12628
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 15304 12628 15332 12656
rect 13872 12600 15332 12628
rect 15473 12631 15531 12637
rect 13872 12588 13878 12600
rect 15473 12597 15485 12631
rect 15519 12628 15531 12631
rect 15562 12628 15568 12640
rect 15519 12600 15568 12628
rect 15519 12597 15531 12600
rect 15473 12591 15531 12597
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 15672 12628 15700 12736
rect 16022 12724 16028 12776
rect 16080 12764 16086 12776
rect 16504 12764 16532 12804
rect 16853 12801 16865 12804
rect 16899 12832 16911 12835
rect 17034 12832 17040 12844
rect 16899 12804 17040 12832
rect 16899 12801 16911 12804
rect 16853 12795 16911 12801
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 17402 12832 17408 12844
rect 17267 12804 17408 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 17880 12841 17908 12872
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 16080 12736 16532 12764
rect 16080 12724 16086 12736
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 17770 12764 17776 12776
rect 16632 12736 17776 12764
rect 16632 12724 16638 12736
rect 17770 12724 17776 12736
rect 17828 12764 17834 12776
rect 17957 12767 18015 12773
rect 17957 12764 17969 12767
rect 17828 12736 17969 12764
rect 17828 12724 17834 12736
rect 17957 12733 17969 12736
rect 18003 12733 18015 12767
rect 17957 12727 18015 12733
rect 15933 12699 15991 12705
rect 15933 12665 15945 12699
rect 15979 12696 15991 12699
rect 15979 12668 16252 12696
rect 15979 12665 15991 12668
rect 15933 12659 15991 12665
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15672 12600 16129 12628
rect 16117 12597 16129 12600
rect 16163 12597 16175 12631
rect 16224 12628 16252 12668
rect 16298 12656 16304 12708
rect 16356 12696 16362 12708
rect 18233 12699 18291 12705
rect 18233 12696 18245 12699
rect 16356 12668 18245 12696
rect 16356 12656 16362 12668
rect 18233 12665 18245 12668
rect 18279 12665 18291 12699
rect 18233 12659 18291 12665
rect 16482 12628 16488 12640
rect 16224 12600 16488 12628
rect 16117 12591 16175 12597
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 17218 12628 17224 12640
rect 17179 12600 17224 12628
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17954 12628 17960 12640
rect 17915 12600 17960 12628
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 1104 12538 18860 12560
rect 1104 12486 3169 12538
rect 3221 12486 3233 12538
rect 3285 12486 3297 12538
rect 3349 12486 3361 12538
rect 3413 12486 3425 12538
rect 3477 12486 7608 12538
rect 7660 12486 7672 12538
rect 7724 12486 7736 12538
rect 7788 12486 7800 12538
rect 7852 12486 7864 12538
rect 7916 12486 12047 12538
rect 12099 12486 12111 12538
rect 12163 12486 12175 12538
rect 12227 12486 12239 12538
rect 12291 12486 12303 12538
rect 12355 12486 16486 12538
rect 16538 12486 16550 12538
rect 16602 12486 16614 12538
rect 16666 12486 16678 12538
rect 16730 12486 16742 12538
rect 16794 12486 18860 12538
rect 1104 12464 18860 12486
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 12345 12427 12403 12433
rect 12345 12424 12357 12427
rect 11388 12396 12357 12424
rect 11388 12384 11394 12396
rect 12345 12393 12357 12396
rect 12391 12424 12403 12427
rect 13814 12424 13820 12436
rect 12391 12396 13820 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 15010 12424 15016 12436
rect 14148 12396 15016 12424
rect 14148 12384 14154 12396
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15654 12384 15660 12436
rect 15712 12424 15718 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 15712 12396 16773 12424
rect 15712 12384 15718 12396
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 17862 12424 17868 12436
rect 16761 12387 16819 12393
rect 17328 12396 17868 12424
rect 17328 12368 17356 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 10502 12316 10508 12368
rect 10560 12356 10566 12368
rect 10560 12328 13216 12356
rect 10560 12316 10566 12328
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 12713 12291 12771 12297
rect 11664 12260 12434 12288
rect 11664 12248 11670 12260
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 11790 12220 11796 12232
rect 11751 12192 11796 12220
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12220 11943 12223
rect 12250 12220 12256 12232
rect 11931 12192 12256 12220
rect 11931 12189 11943 12192
rect 11885 12183 11943 12189
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 12406 12220 12434 12260
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 13078 12288 13084 12300
rect 12759 12260 13084 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 13188 12229 13216 12328
rect 13446 12316 13452 12368
rect 13504 12356 13510 12368
rect 13725 12359 13783 12365
rect 13725 12356 13737 12359
rect 13504 12328 13737 12356
rect 13504 12316 13510 12328
rect 13725 12325 13737 12328
rect 13771 12325 13783 12359
rect 15470 12356 15476 12368
rect 13725 12319 13783 12325
rect 14752 12328 15476 12356
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 13872 12260 14412 12288
rect 13872 12248 13878 12260
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12406 12192 12541 12220
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 13262 12180 13268 12232
rect 13320 12220 13326 12232
rect 13357 12223 13415 12229
rect 13357 12220 13369 12223
rect 13320 12192 13369 12220
rect 13320 12180 13326 12192
rect 13357 12189 13369 12192
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 14182 12220 14188 12232
rect 13587 12192 14188 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 13449 12155 13507 12161
rect 13449 12121 13461 12155
rect 13495 12152 13507 12155
rect 14384 12152 14412 12260
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 14752 12220 14780 12328
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 15749 12359 15807 12365
rect 15749 12325 15761 12359
rect 15795 12325 15807 12359
rect 15749 12319 15807 12325
rect 14826 12248 14832 12300
rect 14884 12248 14890 12300
rect 14918 12248 14924 12300
rect 14976 12288 14982 12300
rect 15102 12288 15108 12300
rect 14976 12260 15108 12288
rect 14976 12248 14982 12260
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 14691 12192 14780 12220
rect 14844 12220 14872 12248
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14844 12192 15025 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 15562 12220 15568 12232
rect 15335 12192 15568 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 15654 12180 15660 12232
rect 15712 12220 15718 12232
rect 15764 12220 15792 12319
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 16853 12359 16911 12365
rect 16853 12356 16865 12359
rect 16448 12328 16865 12356
rect 16448 12316 16454 12328
rect 16853 12325 16865 12328
rect 16899 12325 16911 12359
rect 16853 12319 16911 12325
rect 17310 12316 17316 12368
rect 17368 12316 17374 12368
rect 17586 12316 17592 12368
rect 17644 12356 17650 12368
rect 17773 12359 17831 12365
rect 17773 12356 17785 12359
rect 17644 12328 17785 12356
rect 17644 12316 17650 12328
rect 17773 12325 17785 12328
rect 17819 12325 17831 12359
rect 17773 12319 17831 12325
rect 16114 12288 16120 12300
rect 16040 12260 16120 12288
rect 16040 12229 16068 12260
rect 16114 12248 16120 12260
rect 16172 12248 16178 12300
rect 15712 12192 15792 12220
rect 15933 12223 15991 12229
rect 15712 12180 15718 12192
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16298 12220 16304 12232
rect 16259 12192 16304 12220
rect 16025 12183 16083 12189
rect 14803 12155 14861 12161
rect 14803 12152 14815 12155
rect 13495 12124 13952 12152
rect 14384 12124 14815 12152
rect 13495 12121 13507 12124
rect 13449 12115 13507 12121
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 13814 12084 13820 12096
rect 11296 12056 13820 12084
rect 11296 12044 11302 12056
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 13924 12084 13952 12124
rect 14803 12121 14815 12124
rect 14849 12121 14861 12155
rect 14803 12115 14861 12121
rect 14918 12112 14924 12164
rect 14976 12152 14982 12164
rect 15948 12152 15976 12183
rect 14976 12124 15976 12152
rect 14976 12112 14982 12124
rect 16040 12084 16068 12183
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18138 12220 18144 12232
rect 18003 12192 18144 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 16114 12112 16120 12164
rect 16172 12152 16178 12164
rect 17221 12155 17279 12161
rect 16172 12124 16217 12152
rect 16172 12112 16178 12124
rect 17221 12121 17233 12155
rect 17267 12121 17279 12155
rect 17221 12115 17279 12121
rect 13924 12056 16068 12084
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 17236 12084 17264 12115
rect 16356 12056 17264 12084
rect 16356 12044 16362 12056
rect 1104 11994 19019 12016
rect 1104 11942 5388 11994
rect 5440 11942 5452 11994
rect 5504 11942 5516 11994
rect 5568 11942 5580 11994
rect 5632 11942 5644 11994
rect 5696 11942 9827 11994
rect 9879 11942 9891 11994
rect 9943 11942 9955 11994
rect 10007 11942 10019 11994
rect 10071 11942 10083 11994
rect 10135 11942 14266 11994
rect 14318 11942 14330 11994
rect 14382 11942 14394 11994
rect 14446 11942 14458 11994
rect 14510 11942 14522 11994
rect 14574 11942 18705 11994
rect 18757 11942 18769 11994
rect 18821 11942 18833 11994
rect 18885 11942 18897 11994
rect 18949 11942 18961 11994
rect 19013 11942 19019 11994
rect 1104 11920 19019 11942
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 10928 11852 13093 11880
rect 10928 11840 10934 11852
rect 13081 11849 13093 11852
rect 13127 11849 13139 11883
rect 13906 11880 13912 11892
rect 13867 11852 13912 11880
rect 13081 11843 13139 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 16390 11880 16396 11892
rect 14016 11852 16396 11880
rect 10318 11772 10324 11824
rect 10376 11812 10382 11824
rect 14016 11812 14044 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 18138 11880 18144 11892
rect 18099 11852 18144 11880
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 10376 11784 14044 11812
rect 14185 11815 14243 11821
rect 10376 11772 10382 11784
rect 14185 11781 14197 11815
rect 14231 11781 14243 11815
rect 14185 11775 14243 11781
rect 12618 11744 12624 11756
rect 12579 11716 12624 11744
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 13262 11744 13268 11756
rect 13223 11716 13268 11744
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13372 11716 14105 11744
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 13372 11676 13400 11716
rect 14093 11713 14105 11716
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 10284 11648 13400 11676
rect 13449 11679 13507 11685
rect 10284 11636 10290 11648
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 13814 11676 13820 11688
rect 13495 11648 13820 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 13814 11636 13820 11648
rect 13872 11676 13878 11688
rect 14200 11676 14228 11775
rect 14642 11772 14648 11824
rect 14700 11812 14706 11824
rect 17129 11815 17187 11821
rect 14700 11784 16068 11812
rect 14700 11772 14706 11784
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 14458 11744 14464 11756
rect 14419 11716 14464 11744
rect 14277 11707 14335 11713
rect 13872 11648 14228 11676
rect 13872 11636 13878 11648
rect 10778 11568 10784 11620
rect 10836 11608 10842 11620
rect 14292 11608 14320 11707
rect 14458 11704 14464 11716
rect 14516 11744 14522 11756
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14516 11716 15117 11744
rect 14516 11704 14522 11716
rect 15105 11713 15117 11716
rect 15151 11713 15163 11747
rect 15105 11707 15163 11713
rect 15194 11704 15200 11756
rect 15252 11744 15258 11756
rect 16040 11753 16068 11784
rect 17129 11781 17141 11815
rect 17175 11812 17187 11815
rect 17770 11812 17776 11824
rect 17175 11784 17776 11812
rect 17175 11781 17187 11784
rect 17129 11775 17187 11781
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 15252 11716 15485 11744
rect 15252 11704 15258 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15473 11707 15531 11713
rect 15672 11716 15945 11744
rect 15672 11608 15700 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16908 11716 16957 11744
rect 16908 11704 16914 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 18322 11744 18328 11756
rect 17727 11716 18328 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 10836 11580 14320 11608
rect 14936 11580 15700 11608
rect 10836 11568 10842 11580
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 14936 11549 14964 11580
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 12308 11512 14933 11540
rect 12308 11500 12314 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 15378 11540 15384 11552
rect 15339 11512 15384 11540
rect 14921 11503 14979 11509
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 15933 11543 15991 11549
rect 15933 11540 15945 11543
rect 15804 11512 15945 11540
rect 15804 11500 15810 11512
rect 15933 11509 15945 11512
rect 15979 11509 15991 11543
rect 15933 11503 15991 11509
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16172 11512 16313 11540
rect 16172 11500 16178 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 1104 11450 18860 11472
rect 1104 11398 3169 11450
rect 3221 11398 3233 11450
rect 3285 11398 3297 11450
rect 3349 11398 3361 11450
rect 3413 11398 3425 11450
rect 3477 11398 7608 11450
rect 7660 11398 7672 11450
rect 7724 11398 7736 11450
rect 7788 11398 7800 11450
rect 7852 11398 7864 11450
rect 7916 11398 12047 11450
rect 12099 11398 12111 11450
rect 12163 11398 12175 11450
rect 12227 11398 12239 11450
rect 12291 11398 12303 11450
rect 12355 11398 16486 11450
rect 16538 11398 16550 11450
rect 16602 11398 16614 11450
rect 16666 11398 16678 11450
rect 16730 11398 16742 11450
rect 16794 11398 18860 11450
rect 1104 11376 18860 11398
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 11940 11308 13645 11336
rect 11940 11296 11946 11308
rect 13633 11305 13645 11308
rect 13679 11305 13691 11339
rect 14274 11336 14280 11348
rect 14235 11308 14280 11336
rect 13633 11299 13691 11305
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 15856 11308 16313 11336
rect 14461 11271 14519 11277
rect 14461 11237 14473 11271
rect 14507 11268 14519 11271
rect 15746 11268 15752 11280
rect 14507 11240 15752 11268
rect 14507 11237 14519 11240
rect 14461 11231 14519 11237
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 14476 11200 14504 11231
rect 15746 11228 15752 11240
rect 15804 11228 15810 11280
rect 10468 11172 14504 11200
rect 10468 11160 10474 11172
rect 13556 11141 13584 11172
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14700 11172 14749 11200
rect 14700 11160 14706 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 15856 11200 15884 11308
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 16301 11299 16359 11305
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 17000 11308 17141 11336
rect 17000 11296 17006 11308
rect 17129 11305 17141 11308
rect 17175 11305 17187 11339
rect 18322 11336 18328 11348
rect 18283 11308 18328 11336
rect 17129 11299 17187 11305
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 16132 11240 17172 11268
rect 16132 11209 16160 11240
rect 17144 11212 17172 11240
rect 15068 11172 15884 11200
rect 16117 11203 16175 11209
rect 15068 11160 15074 11172
rect 16117 11169 16129 11203
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 16316 11172 17080 11200
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 13780 11104 13825 11132
rect 13780 11092 13786 11104
rect 15746 11092 15752 11144
rect 15804 11132 15810 11144
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 15804 11104 16221 11132
rect 15804 11092 15810 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 15565 11067 15623 11073
rect 13504 11036 15516 11064
rect 13504 11024 13510 11036
rect 15488 10996 15516 11036
rect 15565 11033 15577 11067
rect 15611 11064 15623 11067
rect 16316 11064 16344 11172
rect 16390 11092 16396 11144
rect 16448 11134 16454 11144
rect 16945 11135 17003 11141
rect 16448 11132 16620 11134
rect 16945 11132 16957 11135
rect 16448 11106 16957 11132
rect 16448 11092 16454 11106
rect 16592 11104 16957 11106
rect 16945 11101 16957 11104
rect 16991 11101 17003 11135
rect 17052 11132 17080 11172
rect 17126 11160 17132 11212
rect 17184 11160 17190 11212
rect 17586 11132 17592 11144
rect 17052 11104 17592 11132
rect 16945 11095 17003 11101
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 16482 11064 16488 11076
rect 15611 11036 16344 11064
rect 16443 11036 16488 11064
rect 15611 11033 15623 11036
rect 15565 11027 15623 11033
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 16114 10996 16120 11008
rect 15488 10968 16120 10996
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 16206 10956 16212 11008
rect 16264 10996 16270 11008
rect 16393 10999 16451 11005
rect 16393 10996 16405 10999
rect 16264 10968 16405 10996
rect 16264 10956 16270 10968
rect 16393 10965 16405 10968
rect 16439 10965 16451 10999
rect 16393 10959 16451 10965
rect 1104 10906 19019 10928
rect 1104 10854 5388 10906
rect 5440 10854 5452 10906
rect 5504 10854 5516 10906
rect 5568 10854 5580 10906
rect 5632 10854 5644 10906
rect 5696 10854 9827 10906
rect 9879 10854 9891 10906
rect 9943 10854 9955 10906
rect 10007 10854 10019 10906
rect 10071 10854 10083 10906
rect 10135 10854 14266 10906
rect 14318 10854 14330 10906
rect 14382 10854 14394 10906
rect 14446 10854 14458 10906
rect 14510 10854 14522 10906
rect 14574 10854 18705 10906
rect 18757 10854 18769 10906
rect 18821 10854 18833 10906
rect 18885 10854 18897 10906
rect 18949 10854 18961 10906
rect 19013 10854 19019 10906
rect 1104 10832 19019 10854
rect 14182 10792 14188 10804
rect 14143 10764 14188 10792
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 15102 10792 15108 10804
rect 15063 10764 15108 10792
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 15565 10795 15623 10801
rect 15565 10761 15577 10795
rect 15611 10792 15623 10795
rect 16850 10792 16856 10804
rect 15611 10764 16856 10792
rect 15611 10761 15623 10764
rect 15565 10755 15623 10761
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17954 10792 17960 10804
rect 16991 10764 17960 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 14826 10724 14832 10736
rect 14752 10696 14832 10724
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14752 10665 14780 10696
rect 14826 10684 14832 10696
rect 14884 10724 14890 10736
rect 16482 10724 16488 10736
rect 14884 10696 16488 10724
rect 14884 10684 14890 10696
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 17126 10724 17132 10736
rect 16868 10696 17132 10724
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 14056 10628 14289 10656
rect 14056 10616 14062 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10625 14795 10659
rect 15838 10656 15844 10668
rect 15799 10628 15844 10656
rect 14737 10619 14795 10625
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16022 10656 16028 10668
rect 15979 10628 16028 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 16868 10665 16896 10696
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17494 10656 17500 10668
rect 17083 10628 17500 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17678 10656 17684 10668
rect 17639 10628 17684 10656
rect 17678 10616 17684 10628
rect 17736 10616 17742 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 18414 10656 18420 10668
rect 18371 10628 18420 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 1578 10588 1584 10600
rect 1539 10560 1584 10588
rect 1578 10548 1584 10560
rect 1636 10548 1642 10600
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 15746 10588 15752 10600
rect 14875 10560 15752 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 14921 10455 14979 10461
rect 14921 10421 14933 10455
rect 14967 10452 14979 10455
rect 15010 10452 15016 10464
rect 14967 10424 15016 10452
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 15933 10455 15991 10461
rect 15933 10421 15945 10455
rect 15979 10452 15991 10455
rect 17218 10452 17224 10464
rect 15979 10424 17224 10452
rect 15979 10421 15991 10424
rect 15933 10415 15991 10421
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 1104 10362 18860 10384
rect 1104 10310 3169 10362
rect 3221 10310 3233 10362
rect 3285 10310 3297 10362
rect 3349 10310 3361 10362
rect 3413 10310 3425 10362
rect 3477 10310 7608 10362
rect 7660 10310 7672 10362
rect 7724 10310 7736 10362
rect 7788 10310 7800 10362
rect 7852 10310 7864 10362
rect 7916 10310 12047 10362
rect 12099 10310 12111 10362
rect 12163 10310 12175 10362
rect 12227 10310 12239 10362
rect 12291 10310 12303 10362
rect 12355 10310 16486 10362
rect 16538 10310 16550 10362
rect 16602 10310 16614 10362
rect 16666 10310 16678 10362
rect 16730 10310 16742 10362
rect 16794 10310 18860 10362
rect 1104 10288 18860 10310
rect 15930 10248 15936 10260
rect 15891 10220 15936 10248
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 17034 10248 17040 10260
rect 16995 10220 17040 10248
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 18322 10248 18328 10260
rect 18283 10220 18328 10248
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 1578 10180 1584 10192
rect 1539 10152 1584 10180
rect 1578 10140 1584 10152
rect 1636 10140 1642 10192
rect 15105 10183 15163 10189
rect 15105 10149 15117 10183
rect 15151 10180 15163 10183
rect 16390 10180 16396 10192
rect 15151 10152 16396 10180
rect 15151 10149 15163 10152
rect 15105 10143 15163 10149
rect 16390 10140 16396 10152
rect 16448 10140 16454 10192
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 14792 10084 15148 10112
rect 14792 10072 14798 10084
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 15120 10053 15148 10084
rect 14921 10047 14979 10053
rect 14921 10044 14933 10047
rect 13688 10016 14933 10044
rect 13688 10004 13694 10016
rect 14921 10013 14933 10016
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 15105 10047 15163 10053
rect 15105 10013 15117 10047
rect 15151 10013 15163 10047
rect 15105 10007 15163 10013
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 17402 10044 17408 10056
rect 17000 10016 17408 10044
rect 17000 10004 17006 10016
rect 17402 10004 17408 10016
rect 17460 10044 17466 10056
rect 17681 10047 17739 10053
rect 17681 10044 17693 10047
rect 17460 10016 17693 10044
rect 17460 10004 17466 10016
rect 17681 10013 17693 10016
rect 17727 10013 17739 10047
rect 17681 10007 17739 10013
rect 1104 9818 19019 9840
rect 1104 9766 5388 9818
rect 5440 9766 5452 9818
rect 5504 9766 5516 9818
rect 5568 9766 5580 9818
rect 5632 9766 5644 9818
rect 5696 9766 9827 9818
rect 9879 9766 9891 9818
rect 9943 9766 9955 9818
rect 10007 9766 10019 9818
rect 10071 9766 10083 9818
rect 10135 9766 14266 9818
rect 14318 9766 14330 9818
rect 14382 9766 14394 9818
rect 14446 9766 14458 9818
rect 14510 9766 14522 9818
rect 14574 9766 18705 9818
rect 18757 9766 18769 9818
rect 18821 9766 18833 9818
rect 18885 9766 18897 9818
rect 18949 9766 18961 9818
rect 19013 9766 19019 9818
rect 1104 9744 19019 9766
rect 19150 9636 19156 9648
rect 16316 9608 19156 9636
rect 16316 9577 16344 9608
rect 19150 9596 19156 9608
rect 19208 9596 19214 9648
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9537 16359 9571
rect 17678 9568 17684 9580
rect 17639 9540 17684 9568
rect 16301 9531 16359 9537
rect 17678 9528 17684 9540
rect 17736 9528 17742 9580
rect 18325 9571 18383 9577
rect 18325 9537 18337 9571
rect 18371 9568 18383 9571
rect 18598 9568 18604 9580
rect 18371 9540 18604 9568
rect 18371 9537 18383 9540
rect 18325 9531 18383 9537
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 15657 9503 15715 9509
rect 15657 9469 15669 9503
rect 15703 9500 15715 9503
rect 16942 9500 16948 9512
rect 15703 9472 16948 9500
rect 15703 9469 15715 9472
rect 15657 9463 15715 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17037 9503 17095 9509
rect 17037 9469 17049 9503
rect 17083 9500 17095 9503
rect 19058 9500 19064 9512
rect 17083 9472 19064 9500
rect 17083 9469 17095 9472
rect 17037 9463 17095 9469
rect 19058 9460 19064 9472
rect 19116 9460 19122 9512
rect 6822 9392 6828 9444
rect 6880 9432 6886 9444
rect 18141 9435 18199 9441
rect 18141 9432 18153 9435
rect 6880 9404 18153 9432
rect 6880 9392 6886 9404
rect 18141 9401 18153 9404
rect 18187 9401 18199 9435
rect 18141 9395 18199 9401
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1104 9274 18860 9296
rect 1104 9222 3169 9274
rect 3221 9222 3233 9274
rect 3285 9222 3297 9274
rect 3349 9222 3361 9274
rect 3413 9222 3425 9274
rect 3477 9222 7608 9274
rect 7660 9222 7672 9274
rect 7724 9222 7736 9274
rect 7788 9222 7800 9274
rect 7852 9222 7864 9274
rect 7916 9222 12047 9274
rect 12099 9222 12111 9274
rect 12163 9222 12175 9274
rect 12227 9222 12239 9274
rect 12291 9222 12303 9274
rect 12355 9222 16486 9274
rect 16538 9222 16550 9274
rect 16602 9222 16614 9274
rect 16666 9222 16678 9274
rect 16730 9222 16742 9274
rect 16794 9222 18860 9274
rect 1104 9200 18860 9222
rect 17681 9163 17739 9169
rect 17681 9129 17693 9163
rect 17727 9160 17739 9163
rect 18230 9160 18236 9172
rect 17727 9132 18236 9160
rect 17727 9129 17739 9132
rect 17681 9123 17739 9129
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 18325 9163 18383 9169
rect 18325 9129 18337 9163
rect 18371 9160 18383 9163
rect 18506 9160 18512 9172
rect 18371 9132 18512 9160
rect 18371 9129 18383 9132
rect 18325 9123 18383 9129
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 16393 9095 16451 9101
rect 16393 9061 16405 9095
rect 16439 9092 16451 9095
rect 19242 9092 19248 9104
rect 16439 9064 19248 9092
rect 16439 9061 16451 9064
rect 16393 9055 16451 9061
rect 19242 9052 19248 9064
rect 19300 9052 19306 9104
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 17034 8956 17040 8968
rect 16995 8928 17040 8956
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 1104 8730 19019 8752
rect 1104 8678 5388 8730
rect 5440 8678 5452 8730
rect 5504 8678 5516 8730
rect 5568 8678 5580 8730
rect 5632 8678 5644 8730
rect 5696 8678 9827 8730
rect 9879 8678 9891 8730
rect 9943 8678 9955 8730
rect 10007 8678 10019 8730
rect 10071 8678 10083 8730
rect 10135 8678 14266 8730
rect 14318 8678 14330 8730
rect 14382 8678 14394 8730
rect 14446 8678 14458 8730
rect 14510 8678 14522 8730
rect 14574 8678 18705 8730
rect 18757 8678 18769 8730
rect 18821 8678 18833 8730
rect 18885 8678 18897 8730
rect 18949 8678 18961 8730
rect 19013 8678 19019 8730
rect 1104 8656 19019 8678
rect 17034 8480 17040 8492
rect 16995 8452 17040 8480
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8480 17739 8483
rect 18046 8480 18052 8492
rect 17727 8452 18052 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18322 8480 18328 8492
rect 18283 8452 18328 8480
rect 18322 8440 18328 8452
rect 18380 8440 18386 8492
rect 1578 8344 1584 8356
rect 1539 8316 1584 8344
rect 1578 8304 1584 8316
rect 1636 8304 1642 8356
rect 1104 8186 18860 8208
rect 1104 8134 3169 8186
rect 3221 8134 3233 8186
rect 3285 8134 3297 8186
rect 3349 8134 3361 8186
rect 3413 8134 3425 8186
rect 3477 8134 7608 8186
rect 7660 8134 7672 8186
rect 7724 8134 7736 8186
rect 7788 8134 7800 8186
rect 7852 8134 7864 8186
rect 7916 8134 12047 8186
rect 12099 8134 12111 8186
rect 12163 8134 12175 8186
rect 12227 8134 12239 8186
rect 12291 8134 12303 8186
rect 12355 8134 16486 8186
rect 16538 8134 16550 8186
rect 16602 8134 16614 8186
rect 16666 8134 16678 8186
rect 16730 8134 16742 8186
rect 16794 8134 18860 8186
rect 1104 8112 18860 8134
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 18598 8072 18604 8084
rect 17727 8044 18604 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 18322 7936 18328 7948
rect 18283 7908 18328 7936
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 1104 7642 19019 7664
rect 1104 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 5644 7642
rect 5696 7590 9827 7642
rect 9879 7590 9891 7642
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7590 10083 7642
rect 10135 7590 14266 7642
rect 14318 7590 14330 7642
rect 14382 7590 14394 7642
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7590 18705 7642
rect 18757 7590 18769 7642
rect 18821 7590 18833 7642
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 18322 7392 18328 7404
rect 18283 7364 18328 7392
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 18322 6780 18328 6792
rect 18283 6752 18328 6780
rect 18322 6740 18328 6752
rect 18380 6740 18386 6792
rect 1104 6554 19019 6576
rect 1104 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 5644 6554
rect 5696 6502 9827 6554
rect 9879 6502 9891 6554
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6502 10083 6554
rect 10135 6502 14266 6554
rect 14318 6502 14330 6554
rect 14382 6502 14394 6554
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6502 18705 6554
rect 18757 6502 18769 6554
rect 18821 6502 18833 6554
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 18322 6304 18328 6316
rect 18283 6276 18328 6304
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 1104 5466 19019 5488
rect 1104 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 5644 5466
rect 5696 5414 9827 5466
rect 9879 5414 9891 5466
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5414 10083 5466
rect 10135 5414 14266 5466
rect 14318 5414 14330 5466
rect 14382 5414 14394 5466
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5414 18705 5466
rect 18757 5414 18769 5466
rect 18821 5414 18833 5466
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 1578 5216 1584 5228
rect 1539 5188 1584 5216
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 18322 5080 18328 5092
rect 18283 5052 18328 5080
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 19150 4604 19156 4616
rect 18371 4576 19156 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 1104 4378 19019 4400
rect 1104 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 5644 4378
rect 5696 4326 9827 4378
rect 9879 4326 9891 4378
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4326 10083 4378
rect 10135 4326 14266 4378
rect 14318 4326 14330 4378
rect 14382 4326 14394 4378
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4326 18705 4378
rect 18757 4326 18769 4378
rect 18821 4326 18833 4378
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 1578 4060 1584 4072
rect 1539 4032 1584 4060
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 18322 3924 18328 3936
rect 18283 3896 18328 3924
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 18322 3516 18328 3528
rect 18283 3488 18328 3516
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 1104 3290 19019 3312
rect 1104 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 5644 3290
rect 5696 3238 9827 3290
rect 9879 3238 9891 3290
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3238 10083 3290
rect 10135 3238 14266 3290
rect 14318 3238 14330 3290
rect 14382 3238 14394 3290
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3238 18705 3290
rect 18757 3238 18769 3290
rect 18821 3238 18833 3290
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 18322 2836 18328 2848
rect 18283 2808 18328 2836
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 2222 2428 2228 2440
rect 2183 2400 2228 2428
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 17678 2428 17684 2440
rect 17639 2400 17684 2428
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 18322 2428 18328 2440
rect 18283 2400 18328 2428
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 1104 2202 19019 2224
rect 1104 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 5644 2202
rect 5696 2150 9827 2202
rect 9879 2150 9891 2202
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2150 10083 2202
rect 10135 2150 14266 2202
rect 14318 2150 14330 2202
rect 14382 2150 14394 2202
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2150 18705 2202
rect 18757 2150 18769 2202
rect 18821 2150 18833 2202
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
<< via1 >>
rect 8116 17824 8168 17876
rect 10416 17824 10468 17876
rect 17132 17824 17184 17876
rect 6184 17756 6236 17808
rect 14648 17756 14700 17808
rect 9404 17688 9456 17740
rect 13728 17688 13780 17740
rect 8484 17552 8536 17604
rect 10232 17552 10284 17604
rect 4712 17484 4764 17536
rect 13636 17484 13688 17536
rect 5388 17382 5440 17434
rect 5452 17382 5504 17434
rect 5516 17382 5568 17434
rect 5580 17382 5632 17434
rect 5644 17382 5696 17434
rect 9827 17382 9879 17434
rect 9891 17382 9943 17434
rect 9955 17382 10007 17434
rect 10019 17382 10071 17434
rect 10083 17382 10135 17434
rect 14266 17382 14318 17434
rect 14330 17382 14382 17434
rect 14394 17382 14446 17434
rect 14458 17382 14510 17434
rect 14522 17382 14574 17434
rect 18705 17382 18757 17434
rect 18769 17382 18821 17434
rect 18833 17382 18885 17434
rect 18897 17382 18949 17434
rect 18961 17382 19013 17434
rect 5724 17280 5776 17332
rect 7564 17280 7616 17332
rect 11796 17280 11848 17332
rect 8116 17212 8168 17264
rect 8300 17212 8352 17264
rect 14188 17280 14240 17332
rect 14280 17280 14332 17332
rect 12992 17212 13044 17264
rect 14740 17212 14792 17264
rect 3332 17144 3384 17196
rect 4804 17144 4856 17196
rect 5172 17144 5224 17196
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 7380 17144 7432 17196
rect 8576 17187 8628 17196
rect 8576 17153 8585 17187
rect 8585 17153 8619 17187
rect 8619 17153 8628 17187
rect 8576 17144 8628 17153
rect 10416 17187 10468 17196
rect 8392 17119 8444 17128
rect 8392 17085 8401 17119
rect 8401 17085 8435 17119
rect 8435 17085 8444 17119
rect 8392 17076 8444 17085
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 11060 17144 11112 17196
rect 13728 17187 13780 17196
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 17040 17212 17092 17264
rect 17224 17212 17276 17264
rect 13728 17144 13780 17153
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 9220 17008 9272 17060
rect 12808 17076 12860 17128
rect 13452 17119 13504 17128
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 14188 17076 14240 17128
rect 16396 17076 16448 17128
rect 1400 16940 1452 16992
rect 6644 16940 6696 16992
rect 7104 16940 7156 16992
rect 8484 16940 8536 16992
rect 9128 16940 9180 16992
rect 11060 17008 11112 17060
rect 17592 17051 17644 17060
rect 9680 16940 9732 16992
rect 10232 16940 10284 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 10876 16940 10928 16992
rect 13728 16940 13780 16992
rect 14648 16940 14700 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 17592 17017 17601 17051
rect 17601 17017 17635 17051
rect 17635 17017 17644 17051
rect 17592 17008 17644 17017
rect 3169 16838 3221 16890
rect 3233 16838 3285 16890
rect 3297 16838 3349 16890
rect 3361 16838 3413 16890
rect 3425 16838 3477 16890
rect 7608 16838 7660 16890
rect 7672 16838 7724 16890
rect 7736 16838 7788 16890
rect 7800 16838 7852 16890
rect 7864 16838 7916 16890
rect 12047 16838 12099 16890
rect 12111 16838 12163 16890
rect 12175 16838 12227 16890
rect 12239 16838 12291 16890
rect 12303 16838 12355 16890
rect 16486 16838 16538 16890
rect 16550 16838 16602 16890
rect 16614 16838 16666 16890
rect 16678 16838 16730 16890
rect 16742 16838 16794 16890
rect 2596 16736 2648 16788
rect 4712 16779 4764 16788
rect 4712 16745 4721 16779
rect 4721 16745 4755 16779
rect 4755 16745 4764 16779
rect 4712 16736 4764 16745
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 8116 16736 8168 16788
rect 8392 16736 8444 16788
rect 10048 16736 10100 16788
rect 10232 16736 10284 16788
rect 10324 16736 10376 16788
rect 13452 16736 13504 16788
rect 13912 16736 13964 16788
rect 16120 16736 16172 16788
rect 6644 16668 6696 16720
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 8300 16532 8352 16584
rect 6000 16507 6052 16516
rect 6000 16473 6009 16507
rect 6009 16473 6043 16507
rect 6043 16473 6052 16507
rect 6000 16464 6052 16473
rect 6644 16507 6696 16516
rect 6644 16473 6653 16507
rect 6653 16473 6687 16507
rect 6687 16473 6696 16507
rect 6644 16464 6696 16473
rect 7840 16464 7892 16516
rect 7104 16396 7156 16448
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 8760 16600 8812 16652
rect 10048 16643 10100 16652
rect 10048 16609 10057 16643
rect 10057 16609 10091 16643
rect 10091 16609 10100 16643
rect 11060 16643 11112 16652
rect 10048 16600 10100 16609
rect 11060 16609 11069 16643
rect 11069 16609 11103 16643
rect 11103 16609 11112 16643
rect 11060 16600 11112 16609
rect 12256 16643 12308 16652
rect 9772 16464 9824 16516
rect 9312 16396 9364 16448
rect 9588 16439 9640 16448
rect 9588 16405 9597 16439
rect 9597 16405 9631 16439
rect 9631 16405 9640 16439
rect 9588 16396 9640 16405
rect 10416 16532 10468 16584
rect 10968 16575 11020 16584
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 10600 16464 10652 16516
rect 11336 16532 11388 16584
rect 10692 16396 10744 16448
rect 11888 16396 11940 16448
rect 12256 16609 12265 16643
rect 12265 16609 12299 16643
rect 12299 16609 12308 16643
rect 12256 16600 12308 16609
rect 12348 16600 12400 16652
rect 14924 16600 14976 16652
rect 16764 16643 16816 16652
rect 13544 16532 13596 16584
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 16764 16609 16773 16643
rect 16773 16609 16807 16643
rect 16807 16609 16816 16643
rect 16764 16600 16816 16609
rect 14004 16464 14056 16516
rect 16120 16532 16172 16584
rect 13176 16396 13228 16448
rect 13544 16396 13596 16448
rect 13820 16396 13872 16448
rect 14740 16396 14792 16448
rect 15476 16396 15528 16448
rect 17316 16464 17368 16516
rect 18328 16464 18380 16516
rect 18236 16439 18288 16448
rect 18236 16405 18245 16439
rect 18245 16405 18279 16439
rect 18279 16405 18288 16439
rect 18236 16396 18288 16405
rect 5388 16294 5440 16346
rect 5452 16294 5504 16346
rect 5516 16294 5568 16346
rect 5580 16294 5632 16346
rect 5644 16294 5696 16346
rect 9827 16294 9879 16346
rect 9891 16294 9943 16346
rect 9955 16294 10007 16346
rect 10019 16294 10071 16346
rect 10083 16294 10135 16346
rect 14266 16294 14318 16346
rect 14330 16294 14382 16346
rect 14394 16294 14446 16346
rect 14458 16294 14510 16346
rect 14522 16294 14574 16346
rect 18705 16294 18757 16346
rect 18769 16294 18821 16346
rect 18833 16294 18885 16346
rect 18897 16294 18949 16346
rect 18961 16294 19013 16346
rect 1124 16056 1176 16108
rect 2872 16099 2924 16108
rect 2872 16065 2881 16099
rect 2881 16065 2915 16099
rect 2915 16065 2924 16099
rect 2872 16056 2924 16065
rect 5172 16099 5224 16108
rect 5172 16065 5181 16099
rect 5181 16065 5215 16099
rect 5215 16065 5224 16099
rect 5172 16056 5224 16065
rect 5356 16099 5408 16108
rect 5356 16065 5365 16099
rect 5365 16065 5399 16099
rect 5399 16065 5408 16099
rect 5356 16056 5408 16065
rect 6828 16167 6880 16176
rect 6828 16133 6855 16167
rect 6855 16133 6880 16167
rect 6828 16124 6880 16133
rect 7104 16124 7156 16176
rect 7196 16124 7248 16176
rect 8576 16192 8628 16244
rect 388 15988 440 16040
rect 6644 15988 6696 16040
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 8300 16056 8352 16108
rect 9956 16124 10008 16176
rect 13268 16192 13320 16244
rect 13820 16192 13872 16244
rect 15844 16192 15896 16244
rect 14924 16124 14976 16176
rect 17040 16167 17092 16176
rect 17040 16133 17049 16167
rect 17049 16133 17083 16167
rect 17083 16133 17092 16167
rect 17040 16124 17092 16133
rect 17592 16167 17644 16176
rect 17592 16133 17601 16167
rect 17601 16133 17635 16167
rect 17635 16133 17644 16167
rect 17592 16124 17644 16133
rect 9036 16056 9088 16108
rect 10784 16056 10836 16108
rect 10968 16056 11020 16108
rect 7840 15988 7892 16040
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8944 16031 8996 16040
rect 8668 15988 8720 15997
rect 8944 15997 8953 16031
rect 8953 15997 8987 16031
rect 8987 15997 8996 16031
rect 8944 15988 8996 15997
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 5264 15852 5316 15904
rect 6000 15895 6052 15904
rect 6000 15861 6009 15895
rect 6009 15861 6043 15895
rect 6043 15861 6052 15895
rect 6000 15852 6052 15861
rect 6736 15852 6788 15904
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 7472 15895 7524 15904
rect 6828 15852 6880 15861
rect 7472 15861 7481 15895
rect 7481 15861 7515 15895
rect 7515 15861 7524 15895
rect 7472 15852 7524 15861
rect 8208 15852 8260 15904
rect 10416 15852 10468 15904
rect 10876 15852 10928 15904
rect 11796 16056 11848 16108
rect 13176 16056 13228 16108
rect 14740 16056 14792 16108
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 11888 15988 11940 16040
rect 14832 15988 14884 16040
rect 15016 15988 15068 16040
rect 15384 15988 15436 16040
rect 14648 15920 14700 15972
rect 12440 15852 12492 15904
rect 12532 15852 12584 15904
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 16304 16031 16356 16040
rect 16304 15997 16313 16031
rect 16313 15997 16347 16031
rect 16347 15997 16356 16031
rect 16304 15988 16356 15997
rect 17224 15988 17276 16040
rect 16396 15920 16448 15972
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 3169 15750 3221 15802
rect 3233 15750 3285 15802
rect 3297 15750 3349 15802
rect 3361 15750 3413 15802
rect 3425 15750 3477 15802
rect 7608 15750 7660 15802
rect 7672 15750 7724 15802
rect 7736 15750 7788 15802
rect 7800 15750 7852 15802
rect 7864 15750 7916 15802
rect 12047 15750 12099 15802
rect 12111 15750 12163 15802
rect 12175 15750 12227 15802
rect 12239 15750 12291 15802
rect 12303 15750 12355 15802
rect 16486 15750 16538 15802
rect 16550 15750 16602 15802
rect 16614 15750 16666 15802
rect 16678 15750 16730 15802
rect 16742 15750 16794 15802
rect 2780 15648 2832 15700
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 6644 15691 6696 15700
rect 6644 15657 6653 15691
rect 6653 15657 6687 15691
rect 6687 15657 6696 15691
rect 6644 15648 6696 15657
rect 6828 15648 6880 15700
rect 7104 15648 7156 15700
rect 7196 15648 7248 15700
rect 8024 15648 8076 15700
rect 11244 15648 11296 15700
rect 12440 15648 12492 15700
rect 15568 15648 15620 15700
rect 5172 15580 5224 15632
rect 7380 15580 7432 15632
rect 8484 15580 8536 15632
rect 8668 15580 8720 15632
rect 9772 15580 9824 15632
rect 11152 15580 11204 15632
rect 11796 15580 11848 15632
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 6736 15512 6788 15564
rect 9220 15512 9272 15564
rect 9680 15512 9732 15564
rect 10784 15512 10836 15564
rect 6736 15376 6788 15428
rect 7104 15444 7156 15496
rect 8024 15444 8076 15496
rect 9404 15444 9456 15496
rect 12992 15512 13044 15564
rect 14556 15512 14608 15564
rect 15016 15512 15068 15564
rect 18328 15512 18380 15564
rect 13820 15444 13872 15496
rect 14832 15444 14884 15496
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 8852 15308 8904 15360
rect 9036 15308 9088 15360
rect 9680 15308 9732 15360
rect 12624 15308 12676 15360
rect 13176 15376 13228 15428
rect 14004 15308 14056 15360
rect 15016 15376 15068 15428
rect 17316 15376 17368 15428
rect 18420 15308 18472 15360
rect 5388 15206 5440 15258
rect 5452 15206 5504 15258
rect 5516 15206 5568 15258
rect 5580 15206 5632 15258
rect 5644 15206 5696 15258
rect 9827 15206 9879 15258
rect 9891 15206 9943 15258
rect 9955 15206 10007 15258
rect 10019 15206 10071 15258
rect 10083 15206 10135 15258
rect 14266 15206 14318 15258
rect 14330 15206 14382 15258
rect 14394 15206 14446 15258
rect 14458 15206 14510 15258
rect 14522 15206 14574 15258
rect 18705 15206 18757 15258
rect 18769 15206 18821 15258
rect 18833 15206 18885 15258
rect 18897 15206 18949 15258
rect 18961 15206 19013 15258
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 11612 15104 11664 15156
rect 12532 15147 12584 15156
rect 12532 15113 12541 15147
rect 12541 15113 12575 15147
rect 12575 15113 12584 15147
rect 12532 15104 12584 15113
rect 12624 15104 12676 15156
rect 12900 15104 12952 15156
rect 1492 14968 1544 15020
rect 7196 15011 7248 15020
rect 7196 14977 7205 15011
rect 7205 14977 7239 15011
rect 7239 14977 7248 15011
rect 7196 14968 7248 14977
rect 8116 15011 8168 15020
rect 8116 14977 8125 15011
rect 8125 14977 8159 15011
rect 8159 14977 8168 15011
rect 8116 14968 8168 14977
rect 8852 15011 8904 15020
rect 6828 14764 6880 14816
rect 8852 14977 8861 15011
rect 8861 14977 8895 15011
rect 8895 14977 8904 15011
rect 8852 14968 8904 14977
rect 10416 14968 10468 15020
rect 10600 14968 10652 15020
rect 9588 14900 9640 14952
rect 10324 14900 10376 14952
rect 10232 14832 10284 14884
rect 10784 14968 10836 15020
rect 12440 15036 12492 15088
rect 13544 15104 13596 15156
rect 13820 15104 13872 15156
rect 11060 14968 11112 15020
rect 14372 15036 14424 15088
rect 14924 15036 14976 15088
rect 15476 15104 15528 15156
rect 17868 15104 17920 15156
rect 17224 15036 17276 15088
rect 17960 15036 18012 15088
rect 15016 14968 15068 15020
rect 17776 14968 17828 15020
rect 18236 15011 18288 15020
rect 18236 14977 18245 15011
rect 18245 14977 18279 15011
rect 18279 14977 18288 15011
rect 18236 14968 18288 14977
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 11704 14900 11756 14952
rect 11888 14943 11940 14952
rect 11888 14909 11897 14943
rect 11897 14909 11931 14943
rect 11931 14909 11940 14943
rect 11888 14900 11940 14909
rect 9036 14764 9088 14816
rect 10048 14764 10100 14816
rect 10784 14764 10836 14816
rect 11152 14807 11204 14816
rect 11152 14773 11161 14807
rect 11161 14773 11195 14807
rect 11195 14773 11204 14807
rect 11152 14764 11204 14773
rect 11520 14832 11572 14884
rect 12992 14900 13044 14952
rect 15292 14832 15344 14884
rect 13084 14764 13136 14816
rect 16120 14900 16172 14952
rect 17040 14900 17092 14952
rect 17132 14943 17184 14952
rect 17132 14909 17141 14943
rect 17141 14909 17175 14943
rect 17175 14909 17184 14943
rect 17500 14943 17552 14952
rect 17132 14900 17184 14909
rect 17500 14909 17509 14943
rect 17509 14909 17543 14943
rect 17543 14909 17552 14943
rect 17500 14900 17552 14909
rect 16396 14832 16448 14884
rect 17684 14764 17736 14816
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 3169 14662 3221 14714
rect 3233 14662 3285 14714
rect 3297 14662 3349 14714
rect 3361 14662 3413 14714
rect 3425 14662 3477 14714
rect 7608 14662 7660 14714
rect 7672 14662 7724 14714
rect 7736 14662 7788 14714
rect 7800 14662 7852 14714
rect 7864 14662 7916 14714
rect 12047 14662 12099 14714
rect 12111 14662 12163 14714
rect 12175 14662 12227 14714
rect 12239 14662 12291 14714
rect 12303 14662 12355 14714
rect 16486 14662 16538 14714
rect 16550 14662 16602 14714
rect 16614 14662 16666 14714
rect 16678 14662 16730 14714
rect 16742 14662 16794 14714
rect 7012 14560 7064 14612
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 10324 14560 10376 14612
rect 11520 14603 11572 14612
rect 11520 14569 11529 14603
rect 11529 14569 11563 14603
rect 11563 14569 11572 14603
rect 11520 14560 11572 14569
rect 11704 14560 11756 14612
rect 15660 14560 15712 14612
rect 8208 14492 8260 14544
rect 10140 14535 10192 14544
rect 10140 14501 10149 14535
rect 10149 14501 10183 14535
rect 10183 14501 10192 14535
rect 10140 14492 10192 14501
rect 11428 14492 11480 14544
rect 10600 14424 10652 14476
rect 11520 14424 11572 14476
rect 11796 14424 11848 14476
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 7196 14288 7248 14340
rect 10048 14288 10100 14340
rect 8300 14220 8352 14272
rect 9588 14263 9640 14272
rect 9588 14229 9597 14263
rect 9597 14229 9631 14263
rect 9631 14229 9640 14263
rect 9588 14220 9640 14229
rect 10784 14356 10836 14408
rect 11060 14356 11112 14408
rect 13452 14424 13504 14476
rect 13912 14424 13964 14476
rect 14648 14424 14700 14476
rect 15016 14424 15068 14476
rect 17408 14424 17460 14476
rect 17776 14424 17828 14476
rect 17960 14424 18012 14476
rect 11244 14288 11296 14340
rect 11428 14288 11480 14340
rect 12992 14288 13044 14340
rect 13912 14288 13964 14340
rect 15292 14288 15344 14340
rect 11704 14220 11756 14272
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 13084 14220 13136 14272
rect 16212 14288 16264 14340
rect 16856 14288 16908 14340
rect 17776 14288 17828 14340
rect 17684 14220 17736 14272
rect 5388 14118 5440 14170
rect 5452 14118 5504 14170
rect 5516 14118 5568 14170
rect 5580 14118 5632 14170
rect 5644 14118 5696 14170
rect 9827 14118 9879 14170
rect 9891 14118 9943 14170
rect 9955 14118 10007 14170
rect 10019 14118 10071 14170
rect 10083 14118 10135 14170
rect 14266 14118 14318 14170
rect 14330 14118 14382 14170
rect 14394 14118 14446 14170
rect 14458 14118 14510 14170
rect 14522 14118 14574 14170
rect 18705 14118 18757 14170
rect 18769 14118 18821 14170
rect 18833 14118 18885 14170
rect 18897 14118 18949 14170
rect 18961 14118 19013 14170
rect 9588 14016 9640 14068
rect 10508 13948 10560 14000
rect 11244 13948 11296 14000
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 9680 13880 9732 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10600 13880 10652 13932
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 12624 14016 12676 14068
rect 12900 14059 12952 14068
rect 12900 14025 12909 14059
rect 12909 14025 12943 14059
rect 12943 14025 12952 14059
rect 12900 14016 12952 14025
rect 13084 14016 13136 14068
rect 11980 13948 12032 14000
rect 12992 13948 13044 14000
rect 12256 13923 12308 13932
rect 12256 13889 12287 13923
rect 12287 13889 12308 13923
rect 12256 13880 12308 13889
rect 12900 13880 12952 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 7288 13812 7340 13864
rect 10324 13812 10376 13864
rect 11244 13812 11296 13864
rect 13544 13948 13596 14000
rect 14924 13948 14976 14000
rect 15108 14016 15160 14068
rect 15200 13948 15252 14000
rect 16028 13991 16080 14000
rect 16028 13957 16063 13991
rect 16063 13957 16080 13991
rect 16028 13948 16080 13957
rect 7472 13744 7524 13796
rect 14004 13812 14056 13864
rect 14648 13812 14700 13864
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 15660 13812 15712 13864
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 15384 13744 15436 13796
rect 17868 13948 17920 14000
rect 17224 13880 17276 13932
rect 17316 13880 17368 13932
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 10324 13676 10376 13728
rect 10508 13676 10560 13728
rect 11244 13676 11296 13728
rect 11796 13676 11848 13728
rect 13360 13676 13412 13728
rect 15108 13719 15160 13728
rect 15108 13685 15117 13719
rect 15117 13685 15151 13719
rect 15151 13685 15160 13719
rect 15108 13676 15160 13685
rect 17040 13676 17092 13728
rect 18420 13744 18472 13796
rect 17960 13719 18012 13728
rect 17960 13685 17969 13719
rect 17969 13685 18003 13719
rect 18003 13685 18012 13719
rect 17960 13676 18012 13685
rect 18052 13676 18104 13728
rect 18236 13676 18288 13728
rect 3169 13574 3221 13626
rect 3233 13574 3285 13626
rect 3297 13574 3349 13626
rect 3361 13574 3413 13626
rect 3425 13574 3477 13626
rect 7608 13574 7660 13626
rect 7672 13574 7724 13626
rect 7736 13574 7788 13626
rect 7800 13574 7852 13626
rect 7864 13574 7916 13626
rect 12047 13574 12099 13626
rect 12111 13574 12163 13626
rect 12175 13574 12227 13626
rect 12239 13574 12291 13626
rect 12303 13574 12355 13626
rect 16486 13574 16538 13626
rect 16550 13574 16602 13626
rect 16614 13574 16666 13626
rect 16678 13574 16730 13626
rect 16742 13574 16794 13626
rect 11060 13472 11112 13524
rect 6736 13336 6788 13388
rect 10508 13404 10560 13456
rect 11244 13404 11296 13456
rect 11612 13404 11664 13456
rect 11980 13404 12032 13456
rect 12164 13472 12216 13524
rect 16028 13472 16080 13524
rect 17040 13515 17092 13524
rect 17040 13481 17049 13515
rect 17049 13481 17083 13515
rect 17083 13481 17092 13515
rect 17040 13472 17092 13481
rect 17500 13472 17552 13524
rect 17868 13515 17920 13524
rect 17868 13481 17877 13515
rect 17877 13481 17911 13515
rect 17911 13481 17920 13515
rect 17868 13472 17920 13481
rect 12532 13404 12584 13456
rect 13728 13404 13780 13456
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 7104 13268 7156 13320
rect 9864 13268 9916 13320
rect 10600 13268 10652 13320
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 11244 13268 11296 13320
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 11888 13268 11940 13320
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 13176 13336 13228 13388
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13360 13336 13412 13345
rect 13452 13336 13504 13388
rect 16304 13336 16356 13388
rect 16396 13336 16448 13388
rect 13544 13268 13596 13320
rect 13820 13268 13872 13320
rect 15844 13268 15896 13320
rect 17316 13336 17368 13388
rect 17500 13336 17552 13388
rect 16672 13311 16724 13320
rect 12348 13200 12400 13252
rect 15292 13200 15344 13252
rect 8392 13132 8444 13184
rect 10416 13132 10468 13184
rect 11888 13132 11940 13184
rect 11980 13132 12032 13184
rect 12440 13132 12492 13184
rect 12900 13132 12952 13184
rect 16212 13200 16264 13252
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 16396 13200 16448 13252
rect 17132 13243 17184 13252
rect 17132 13209 17141 13243
rect 17141 13209 17175 13243
rect 17175 13209 17184 13243
rect 17132 13200 17184 13209
rect 17684 13200 17736 13252
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 17040 13132 17092 13184
rect 17868 13132 17920 13184
rect 5388 13030 5440 13082
rect 5452 13030 5504 13082
rect 5516 13030 5568 13082
rect 5580 13030 5632 13082
rect 5644 13030 5696 13082
rect 9827 13030 9879 13082
rect 9891 13030 9943 13082
rect 9955 13030 10007 13082
rect 10019 13030 10071 13082
rect 10083 13030 10135 13082
rect 14266 13030 14318 13082
rect 14330 13030 14382 13082
rect 14394 13030 14446 13082
rect 14458 13030 14510 13082
rect 14522 13030 14574 13082
rect 18705 13030 18757 13082
rect 18769 13030 18821 13082
rect 18833 13030 18885 13082
rect 18897 13030 18949 13082
rect 18961 13030 19013 13082
rect 9312 12928 9364 12980
rect 11152 12928 11204 12980
rect 12716 12928 12768 12980
rect 13268 12928 13320 12980
rect 14188 12928 14240 12980
rect 14924 12928 14976 12980
rect 17408 12971 17460 12980
rect 6000 12860 6052 12912
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 11888 12860 11940 12912
rect 15292 12860 15344 12912
rect 16304 12903 16356 12912
rect 16304 12869 16313 12903
rect 16313 12869 16347 12903
rect 16347 12869 16356 12903
rect 16304 12860 16356 12869
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 11060 12792 11112 12844
rect 9036 12656 9088 12708
rect 10968 12699 11020 12708
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 8484 12588 8536 12640
rect 10508 12588 10560 12640
rect 10968 12665 10977 12699
rect 10977 12665 11011 12699
rect 11011 12665 11020 12699
rect 10968 12656 11020 12665
rect 11704 12792 11756 12844
rect 12440 12792 12492 12844
rect 12532 12792 12584 12844
rect 13084 12792 13136 12844
rect 15384 12792 15436 12844
rect 15568 12792 15620 12844
rect 16396 12792 16448 12844
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 11520 12656 11572 12708
rect 12624 12656 12676 12708
rect 15292 12656 15344 12708
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 13820 12588 13872 12640
rect 15568 12588 15620 12640
rect 16028 12724 16080 12776
rect 17040 12792 17092 12844
rect 17408 12792 17460 12844
rect 16580 12724 16632 12776
rect 17776 12724 17828 12776
rect 16304 12656 16356 12708
rect 16488 12588 16540 12640
rect 17224 12631 17276 12640
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 17224 12588 17276 12597
rect 17960 12631 18012 12640
rect 17960 12597 17969 12631
rect 17969 12597 18003 12631
rect 18003 12597 18012 12631
rect 17960 12588 18012 12597
rect 3169 12486 3221 12538
rect 3233 12486 3285 12538
rect 3297 12486 3349 12538
rect 3361 12486 3413 12538
rect 3425 12486 3477 12538
rect 7608 12486 7660 12538
rect 7672 12486 7724 12538
rect 7736 12486 7788 12538
rect 7800 12486 7852 12538
rect 7864 12486 7916 12538
rect 12047 12486 12099 12538
rect 12111 12486 12163 12538
rect 12175 12486 12227 12538
rect 12239 12486 12291 12538
rect 12303 12486 12355 12538
rect 16486 12486 16538 12538
rect 16550 12486 16602 12538
rect 16614 12486 16666 12538
rect 16678 12486 16730 12538
rect 16742 12486 16794 12538
rect 11336 12384 11388 12436
rect 13820 12384 13872 12436
rect 14096 12384 14148 12436
rect 15016 12427 15068 12436
rect 15016 12393 15025 12427
rect 15025 12393 15059 12427
rect 15059 12393 15068 12427
rect 15016 12384 15068 12393
rect 15660 12384 15712 12436
rect 17868 12384 17920 12436
rect 10508 12316 10560 12368
rect 11612 12248 11664 12300
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 12256 12180 12308 12232
rect 13084 12248 13136 12300
rect 13452 12316 13504 12368
rect 13820 12248 13872 12300
rect 13268 12180 13320 12232
rect 14188 12180 14240 12232
rect 15476 12316 15528 12368
rect 14832 12248 14884 12300
rect 14924 12248 14976 12300
rect 15108 12248 15160 12300
rect 15568 12180 15620 12232
rect 15660 12180 15712 12232
rect 16396 12316 16448 12368
rect 17316 12316 17368 12368
rect 17592 12316 17644 12368
rect 16120 12248 16172 12300
rect 16304 12223 16356 12232
rect 11244 12044 11296 12096
rect 13820 12044 13872 12096
rect 14924 12112 14976 12164
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 18144 12180 18196 12232
rect 16120 12155 16172 12164
rect 16120 12121 16129 12155
rect 16129 12121 16163 12155
rect 16163 12121 16172 12155
rect 16120 12112 16172 12121
rect 16304 12044 16356 12096
rect 5388 11942 5440 11994
rect 5452 11942 5504 11994
rect 5516 11942 5568 11994
rect 5580 11942 5632 11994
rect 5644 11942 5696 11994
rect 9827 11942 9879 11994
rect 9891 11942 9943 11994
rect 9955 11942 10007 11994
rect 10019 11942 10071 11994
rect 10083 11942 10135 11994
rect 14266 11942 14318 11994
rect 14330 11942 14382 11994
rect 14394 11942 14446 11994
rect 14458 11942 14510 11994
rect 14522 11942 14574 11994
rect 18705 11942 18757 11994
rect 18769 11942 18821 11994
rect 18833 11942 18885 11994
rect 18897 11942 18949 11994
rect 18961 11942 19013 11994
rect 10876 11840 10928 11892
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 10324 11772 10376 11824
rect 16396 11840 16448 11892
rect 18144 11883 18196 11892
rect 18144 11849 18153 11883
rect 18153 11849 18187 11883
rect 18187 11849 18196 11883
rect 18144 11840 18196 11849
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 13268 11747 13320 11756
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 10232 11636 10284 11688
rect 13820 11636 13872 11688
rect 14648 11772 14700 11824
rect 14464 11747 14516 11756
rect 10784 11568 10836 11620
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 15200 11704 15252 11756
rect 17776 11772 17828 11824
rect 16856 11704 16908 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 12256 11500 12308 11552
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 15752 11500 15804 11552
rect 16120 11500 16172 11552
rect 3169 11398 3221 11450
rect 3233 11398 3285 11450
rect 3297 11398 3349 11450
rect 3361 11398 3413 11450
rect 3425 11398 3477 11450
rect 7608 11398 7660 11450
rect 7672 11398 7724 11450
rect 7736 11398 7788 11450
rect 7800 11398 7852 11450
rect 7864 11398 7916 11450
rect 12047 11398 12099 11450
rect 12111 11398 12163 11450
rect 12175 11398 12227 11450
rect 12239 11398 12291 11450
rect 12303 11398 12355 11450
rect 16486 11398 16538 11450
rect 16550 11398 16602 11450
rect 16614 11398 16666 11450
rect 16678 11398 16730 11450
rect 16742 11398 16794 11450
rect 11888 11296 11940 11348
rect 14280 11339 14332 11348
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 10416 11160 10468 11212
rect 15752 11228 15804 11280
rect 14648 11160 14700 11212
rect 15016 11160 15068 11212
rect 16948 11296 17000 11348
rect 18328 11339 18380 11348
rect 18328 11305 18337 11339
rect 18337 11305 18371 11339
rect 18371 11305 18380 11339
rect 18328 11296 18380 11305
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 15752 11092 15804 11144
rect 13452 11024 13504 11076
rect 16396 11092 16448 11144
rect 17132 11160 17184 11212
rect 17592 11092 17644 11144
rect 16488 11067 16540 11076
rect 16488 11033 16497 11067
rect 16497 11033 16531 11067
rect 16531 11033 16540 11067
rect 16488 11024 16540 11033
rect 16120 10956 16172 11008
rect 16212 10956 16264 11008
rect 5388 10854 5440 10906
rect 5452 10854 5504 10906
rect 5516 10854 5568 10906
rect 5580 10854 5632 10906
rect 5644 10854 5696 10906
rect 9827 10854 9879 10906
rect 9891 10854 9943 10906
rect 9955 10854 10007 10906
rect 10019 10854 10071 10906
rect 10083 10854 10135 10906
rect 14266 10854 14318 10906
rect 14330 10854 14382 10906
rect 14394 10854 14446 10906
rect 14458 10854 14510 10906
rect 14522 10854 14574 10906
rect 18705 10854 18757 10906
rect 18769 10854 18821 10906
rect 18833 10854 18885 10906
rect 18897 10854 18949 10906
rect 18961 10854 19013 10906
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 15108 10795 15160 10804
rect 15108 10761 15117 10795
rect 15117 10761 15151 10795
rect 15151 10761 15160 10795
rect 15108 10752 15160 10761
rect 16856 10752 16908 10804
rect 17960 10752 18012 10804
rect 14004 10616 14056 10668
rect 14832 10684 14884 10736
rect 16488 10684 16540 10736
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 16028 10616 16080 10668
rect 17132 10684 17184 10736
rect 17500 10616 17552 10668
rect 17684 10659 17736 10668
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 18420 10616 18472 10668
rect 1584 10591 1636 10600
rect 1584 10557 1593 10591
rect 1593 10557 1627 10591
rect 1627 10557 1636 10591
rect 1584 10548 1636 10557
rect 15752 10548 15804 10600
rect 15016 10412 15068 10464
rect 17224 10412 17276 10464
rect 3169 10310 3221 10362
rect 3233 10310 3285 10362
rect 3297 10310 3349 10362
rect 3361 10310 3413 10362
rect 3425 10310 3477 10362
rect 7608 10310 7660 10362
rect 7672 10310 7724 10362
rect 7736 10310 7788 10362
rect 7800 10310 7852 10362
rect 7864 10310 7916 10362
rect 12047 10310 12099 10362
rect 12111 10310 12163 10362
rect 12175 10310 12227 10362
rect 12239 10310 12291 10362
rect 12303 10310 12355 10362
rect 16486 10310 16538 10362
rect 16550 10310 16602 10362
rect 16614 10310 16666 10362
rect 16678 10310 16730 10362
rect 16742 10310 16794 10362
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 17040 10251 17092 10260
rect 17040 10217 17049 10251
rect 17049 10217 17083 10251
rect 17083 10217 17092 10251
rect 17040 10208 17092 10217
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 1584 10183 1636 10192
rect 1584 10149 1593 10183
rect 1593 10149 1627 10183
rect 1627 10149 1636 10183
rect 1584 10140 1636 10149
rect 16396 10140 16448 10192
rect 14740 10072 14792 10124
rect 13636 10004 13688 10056
rect 16948 10004 17000 10056
rect 17408 10004 17460 10056
rect 5388 9766 5440 9818
rect 5452 9766 5504 9818
rect 5516 9766 5568 9818
rect 5580 9766 5632 9818
rect 5644 9766 5696 9818
rect 9827 9766 9879 9818
rect 9891 9766 9943 9818
rect 9955 9766 10007 9818
rect 10019 9766 10071 9818
rect 10083 9766 10135 9818
rect 14266 9766 14318 9818
rect 14330 9766 14382 9818
rect 14394 9766 14446 9818
rect 14458 9766 14510 9818
rect 14522 9766 14574 9818
rect 18705 9766 18757 9818
rect 18769 9766 18821 9818
rect 18833 9766 18885 9818
rect 18897 9766 18949 9818
rect 18961 9766 19013 9818
rect 19156 9596 19208 9648
rect 17684 9571 17736 9580
rect 17684 9537 17693 9571
rect 17693 9537 17727 9571
rect 17727 9537 17736 9571
rect 17684 9528 17736 9537
rect 18604 9528 18656 9580
rect 16948 9460 17000 9512
rect 19064 9460 19116 9512
rect 6828 9392 6880 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3169 9222 3221 9274
rect 3233 9222 3285 9274
rect 3297 9222 3349 9274
rect 3361 9222 3413 9274
rect 3425 9222 3477 9274
rect 7608 9222 7660 9274
rect 7672 9222 7724 9274
rect 7736 9222 7788 9274
rect 7800 9222 7852 9274
rect 7864 9222 7916 9274
rect 12047 9222 12099 9274
rect 12111 9222 12163 9274
rect 12175 9222 12227 9274
rect 12239 9222 12291 9274
rect 12303 9222 12355 9274
rect 16486 9222 16538 9274
rect 16550 9222 16602 9274
rect 16614 9222 16666 9274
rect 16678 9222 16730 9274
rect 16742 9222 16794 9274
rect 18236 9120 18288 9172
rect 18512 9120 18564 9172
rect 19248 9052 19300 9104
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 17040 8959 17092 8968
rect 17040 8925 17049 8959
rect 17049 8925 17083 8959
rect 17083 8925 17092 8959
rect 17040 8916 17092 8925
rect 5388 8678 5440 8730
rect 5452 8678 5504 8730
rect 5516 8678 5568 8730
rect 5580 8678 5632 8730
rect 5644 8678 5696 8730
rect 9827 8678 9879 8730
rect 9891 8678 9943 8730
rect 9955 8678 10007 8730
rect 10019 8678 10071 8730
rect 10083 8678 10135 8730
rect 14266 8678 14318 8730
rect 14330 8678 14382 8730
rect 14394 8678 14446 8730
rect 14458 8678 14510 8730
rect 14522 8678 14574 8730
rect 18705 8678 18757 8730
rect 18769 8678 18821 8730
rect 18833 8678 18885 8730
rect 18897 8678 18949 8730
rect 18961 8678 19013 8730
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 18052 8440 18104 8492
rect 18328 8483 18380 8492
rect 18328 8449 18337 8483
rect 18337 8449 18371 8483
rect 18371 8449 18380 8483
rect 18328 8440 18380 8449
rect 1584 8347 1636 8356
rect 1584 8313 1593 8347
rect 1593 8313 1627 8347
rect 1627 8313 1636 8347
rect 1584 8304 1636 8313
rect 3169 8134 3221 8186
rect 3233 8134 3285 8186
rect 3297 8134 3349 8186
rect 3361 8134 3413 8186
rect 3425 8134 3477 8186
rect 7608 8134 7660 8186
rect 7672 8134 7724 8186
rect 7736 8134 7788 8186
rect 7800 8134 7852 8186
rect 7864 8134 7916 8186
rect 12047 8134 12099 8186
rect 12111 8134 12163 8186
rect 12175 8134 12227 8186
rect 12239 8134 12291 8186
rect 12303 8134 12355 8186
rect 16486 8134 16538 8186
rect 16550 8134 16602 8186
rect 16614 8134 16666 8186
rect 16678 8134 16730 8186
rect 16742 8134 16794 8186
rect 18604 8032 18656 8084
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 5644 7590 5696 7642
rect 9827 7590 9879 7642
rect 9891 7590 9943 7642
rect 9955 7590 10007 7642
rect 10019 7590 10071 7642
rect 10083 7590 10135 7642
rect 14266 7590 14318 7642
rect 14330 7590 14382 7642
rect 14394 7590 14446 7642
rect 14458 7590 14510 7642
rect 14522 7590 14574 7642
rect 18705 7590 18757 7642
rect 18769 7590 18821 7642
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 18328 6783 18380 6792
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 5644 6502 5696 6554
rect 9827 6502 9879 6554
rect 9891 6502 9943 6554
rect 9955 6502 10007 6554
rect 10019 6502 10071 6554
rect 10083 6502 10135 6554
rect 14266 6502 14318 6554
rect 14330 6502 14382 6554
rect 14394 6502 14446 6554
rect 14458 6502 14510 6554
rect 14522 6502 14574 6554
rect 18705 6502 18757 6554
rect 18769 6502 18821 6554
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 18328 6307 18380 6316
rect 18328 6273 18337 6307
rect 18337 6273 18371 6307
rect 18371 6273 18380 6307
rect 18328 6264 18380 6273
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 5644 5414 5696 5466
rect 9827 5414 9879 5466
rect 9891 5414 9943 5466
rect 9955 5414 10007 5466
rect 10019 5414 10071 5466
rect 10083 5414 10135 5466
rect 14266 5414 14318 5466
rect 14330 5414 14382 5466
rect 14394 5414 14446 5466
rect 14458 5414 14510 5466
rect 14522 5414 14574 5466
rect 18705 5414 18757 5466
rect 18769 5414 18821 5466
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 18328 5083 18380 5092
rect 18328 5049 18337 5083
rect 18337 5049 18371 5083
rect 18371 5049 18380 5083
rect 18328 5040 18380 5049
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 19156 4564 19208 4616
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 5644 4326 5696 4378
rect 9827 4326 9879 4378
rect 9891 4326 9943 4378
rect 9955 4326 10007 4378
rect 10019 4326 10071 4378
rect 10083 4326 10135 4378
rect 14266 4326 14318 4378
rect 14330 4326 14382 4378
rect 14394 4326 14446 4378
rect 14458 4326 14510 4378
rect 14522 4326 14574 4378
rect 18705 4326 18757 4378
rect 18769 4326 18821 4378
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 1584 4063 1636 4072
rect 1584 4029 1593 4063
rect 1593 4029 1627 4063
rect 1627 4029 1636 4063
rect 1584 4020 1636 4029
rect 18328 3927 18380 3936
rect 18328 3893 18337 3927
rect 18337 3893 18371 3927
rect 18371 3893 18380 3927
rect 18328 3884 18380 3893
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 5644 3238 5696 3290
rect 9827 3238 9879 3290
rect 9891 3238 9943 3290
rect 9955 3238 10007 3290
rect 10019 3238 10071 3290
rect 10083 3238 10135 3290
rect 14266 3238 14318 3290
rect 14330 3238 14382 3290
rect 14394 3238 14446 3290
rect 14458 3238 14510 3290
rect 14522 3238 14574 3290
rect 18705 3238 18757 3290
rect 18769 3238 18821 3290
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 5644 2150 5696 2202
rect 9827 2150 9879 2202
rect 9891 2150 9943 2202
rect 9955 2150 10007 2202
rect 10019 2150 10071 2202
rect 10083 2150 10135 2202
rect 14266 2150 14318 2202
rect 14330 2150 14382 2202
rect 14394 2150 14446 2202
rect 14458 2150 14510 2202
rect 14522 2150 14574 2202
rect 18705 2150 18757 2202
rect 18769 2150 18821 2202
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
<< metal2 >>
rect 386 19200 442 20000
rect 1122 19200 1178 20000
rect 1858 19200 1914 20000
rect 2594 19200 2650 20000
rect 3330 19200 3386 20000
rect 4066 19200 4122 20000
rect 4802 19200 4858 20000
rect 5538 19200 5594 20000
rect 6274 19200 6330 20000
rect 7010 19200 7066 20000
rect 7746 19200 7802 20000
rect 8482 19200 8538 20000
rect 9218 19200 9274 20000
rect 9692 19230 9904 19258
rect 400 16046 428 19200
rect 1136 16114 1164 19200
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16697 1440 16934
rect 2608 16794 2636 19200
rect 2778 17912 2834 17921
rect 2778 17847 2834 17856
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 1398 16688 1454 16697
rect 1398 16623 1454 16632
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 16289 1624 16594
rect 1582 16280 1638 16289
rect 1582 16215 1638 16224
rect 1124 16108 1176 16114
rect 1124 16050 1176 16056
rect 388 16040 440 16046
rect 388 15982 440 15988
rect 2792 15706 2820 17847
rect 2870 17504 2926 17513
rect 2870 17439 2926 17448
rect 2884 16114 2912 17439
rect 3344 17202 3372 19200
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3169 16892 3477 16901
rect 3169 16890 3175 16892
rect 3231 16890 3255 16892
rect 3311 16890 3335 16892
rect 3391 16890 3415 16892
rect 3471 16890 3477 16892
rect 3231 16838 3233 16890
rect 3413 16838 3415 16890
rect 3169 16836 3175 16838
rect 3231 16836 3255 16838
rect 3311 16836 3335 16838
rect 3391 16836 3415 16838
rect 3471 16836 3477 16838
rect 3169 16827 3477 16836
rect 4724 16794 4752 17478
rect 4816 17202 4844 19200
rect 5552 17626 5580 19200
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 5552 17598 5764 17626
rect 5388 17436 5696 17445
rect 5388 17434 5394 17436
rect 5450 17434 5474 17436
rect 5530 17434 5554 17436
rect 5610 17434 5634 17436
rect 5690 17434 5696 17436
rect 5450 17382 5452 17434
rect 5632 17382 5634 17434
rect 5388 17380 5394 17382
rect 5450 17380 5474 17382
rect 5530 17380 5554 17382
rect 5610 17380 5634 17382
rect 5690 17380 5696 17382
rect 5388 17371 5696 17380
rect 5736 17338 5764 17598
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 5184 16590 5212 17138
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5998 16552 6054 16561
rect 5998 16487 6000 16496
rect 6052 16487 6054 16496
rect 6000 16458 6052 16464
rect 5388 16348 5696 16357
rect 5388 16346 5394 16348
rect 5450 16346 5474 16348
rect 5530 16346 5554 16348
rect 5610 16346 5634 16348
rect 5690 16346 5696 16348
rect 5450 16294 5452 16346
rect 5632 16294 5634 16346
rect 5388 16292 5394 16294
rect 5450 16292 5474 16294
rect 5530 16292 5554 16294
rect 5610 16292 5634 16294
rect 5690 16292 5696 16294
rect 5388 16283 5696 16292
rect 5354 16144 5410 16153
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 5172 16108 5224 16114
rect 5354 16079 5356 16088
rect 5172 16050 5224 16056
rect 5408 16079 5410 16088
rect 5356 16050 5408 16056
rect 3169 15804 3477 15813
rect 3169 15802 3175 15804
rect 3231 15802 3255 15804
rect 3311 15802 3335 15804
rect 3391 15802 3415 15804
rect 3471 15802 3477 15804
rect 3231 15750 3233 15802
rect 3413 15750 3415 15802
rect 3169 15748 3175 15750
rect 3231 15748 3255 15750
rect 3311 15748 3335 15750
rect 3391 15748 3415 15750
rect 3471 15748 3477 15750
rect 3169 15739 3477 15748
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 5184 15638 5212 16050
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 1584 15496 1636 15502
rect 1490 15464 1546 15473
rect 1584 15438 1636 15444
rect 1490 15399 1546 15408
rect 1504 15026 1532 15399
rect 1596 15065 1624 15438
rect 1582 15056 1638 15065
rect 1492 15020 1544 15026
rect 1582 14991 1638 15000
rect 1492 14962 1544 14968
rect 3169 14716 3477 14725
rect 3169 14714 3175 14716
rect 3231 14714 3255 14716
rect 3311 14714 3335 14716
rect 3391 14714 3415 14716
rect 3471 14714 3477 14716
rect 3231 14662 3233 14714
rect 3413 14662 3415 14714
rect 3169 14660 3175 14662
rect 3231 14660 3255 14662
rect 3311 14660 3335 14662
rect 3391 14660 3415 14662
rect 3471 14660 3477 14662
rect 3169 14651 3477 14660
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 14249 1624 14350
rect 1582 14240 1638 14249
rect 1582 14175 1638 14184
rect 1584 13864 1636 13870
rect 1582 13832 1584 13841
rect 1636 13832 1638 13841
rect 1582 13767 1638 13776
rect 3169 13628 3477 13637
rect 3169 13626 3175 13628
rect 3231 13626 3255 13628
rect 3311 13626 3335 13628
rect 3391 13626 3415 13628
rect 3471 13626 3477 13628
rect 3231 13574 3233 13626
rect 3413 13574 3415 13626
rect 3169 13572 3175 13574
rect 3231 13572 3255 13574
rect 3311 13572 3335 13574
rect 3391 13572 3415 13574
rect 3471 13572 3477 13574
rect 3169 13563 3477 13572
rect 5276 13433 5304 15846
rect 5388 15260 5696 15269
rect 5388 15258 5394 15260
rect 5450 15258 5474 15260
rect 5530 15258 5554 15260
rect 5610 15258 5634 15260
rect 5690 15258 5696 15260
rect 5450 15206 5452 15258
rect 5632 15206 5634 15258
rect 5388 15204 5394 15206
rect 5450 15204 5474 15206
rect 5530 15204 5554 15206
rect 5610 15204 5634 15206
rect 5690 15204 5696 15206
rect 5388 15195 5696 15204
rect 5388 14172 5696 14181
rect 5388 14170 5394 14172
rect 5450 14170 5474 14172
rect 5530 14170 5554 14172
rect 5610 14170 5634 14172
rect 5690 14170 5696 14172
rect 5450 14118 5452 14170
rect 5632 14118 5634 14170
rect 5388 14116 5394 14118
rect 5450 14116 5474 14118
rect 5530 14116 5554 14118
rect 5610 14116 5634 14118
rect 5690 14116 5696 14118
rect 5388 14107 5696 14116
rect 5262 13424 5318 13433
rect 5262 13359 5318 13368
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 13025 1624 13262
rect 5388 13084 5696 13093
rect 5388 13082 5394 13084
rect 5450 13082 5474 13084
rect 5530 13082 5554 13084
rect 5610 13082 5634 13084
rect 5690 13082 5696 13084
rect 5450 13030 5452 13082
rect 5632 13030 5634 13082
rect 5388 13028 5394 13030
rect 5450 13028 5474 13030
rect 5530 13028 5554 13030
rect 5610 13028 5634 13030
rect 5690 13028 5696 13030
rect 1582 13016 1638 13025
rect 5388 13019 5696 13028
rect 1582 12951 1638 12960
rect 6012 12918 6040 15846
rect 6196 15706 6224 17750
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6656 16726 6684 16934
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6656 16522 6684 16662
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6644 16040 6696 16046
rect 6840 16017 6868 16118
rect 6644 15982 6696 15988
rect 6826 16008 6882 16017
rect 6656 15706 6684 15982
rect 6826 15943 6882 15952
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6748 15570 6776 15846
rect 6840 15706 6868 15846
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6748 13394 6776 15370
rect 6932 14906 6960 17138
rect 6840 14878 6960 14906
rect 6840 14822 6868 14878
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6000 12912 6052 12918
rect 6000 12854 6052 12860
rect 1584 12640 1636 12646
rect 1582 12608 1584 12617
rect 1636 12608 1638 12617
rect 1582 12543 1638 12552
rect 3169 12540 3477 12549
rect 3169 12538 3175 12540
rect 3231 12538 3255 12540
rect 3311 12538 3335 12540
rect 3391 12538 3415 12540
rect 3471 12538 3477 12540
rect 3231 12486 3233 12538
rect 3413 12486 3415 12538
rect 3169 12484 3175 12486
rect 3231 12484 3255 12486
rect 3311 12484 3335 12486
rect 3391 12484 3415 12486
rect 3471 12484 3477 12486
rect 3169 12475 3477 12484
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11801 1624 12174
rect 5388 11996 5696 12005
rect 5388 11994 5394 11996
rect 5450 11994 5474 11996
rect 5530 11994 5554 11996
rect 5610 11994 5634 11996
rect 5690 11994 5696 11996
rect 5450 11942 5452 11994
rect 5632 11942 5634 11994
rect 5388 11940 5394 11942
rect 5450 11940 5474 11942
rect 5530 11940 5554 11942
rect 5610 11940 5634 11942
rect 5690 11940 5696 11942
rect 5388 11931 5696 11940
rect 1582 11792 1638 11801
rect 1582 11727 1638 11736
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11393 1624 11494
rect 3169 11452 3477 11461
rect 3169 11450 3175 11452
rect 3231 11450 3255 11452
rect 3311 11450 3335 11452
rect 3391 11450 3415 11452
rect 3471 11450 3477 11452
rect 3231 11398 3233 11450
rect 3413 11398 3415 11450
rect 3169 11396 3175 11398
rect 3231 11396 3255 11398
rect 3311 11396 3335 11398
rect 3391 11396 3415 11398
rect 3471 11396 3477 11398
rect 1582 11384 1638 11393
rect 3169 11387 3477 11396
rect 1582 11319 1638 11328
rect 5388 10908 5696 10917
rect 5388 10906 5394 10908
rect 5450 10906 5474 10908
rect 5530 10906 5554 10908
rect 5610 10906 5634 10908
rect 5690 10906 5696 10908
rect 5450 10854 5452 10906
rect 5632 10854 5634 10906
rect 5388 10852 5394 10854
rect 5450 10852 5474 10854
rect 5530 10852 5554 10854
rect 5610 10852 5634 10854
rect 5690 10852 5696 10854
rect 5388 10843 5696 10852
rect 1584 10600 1636 10606
rect 1582 10568 1584 10577
rect 1636 10568 1638 10577
rect 1582 10503 1638 10512
rect 3169 10364 3477 10373
rect 3169 10362 3175 10364
rect 3231 10362 3255 10364
rect 3311 10362 3335 10364
rect 3391 10362 3415 10364
rect 3471 10362 3477 10364
rect 3231 10310 3233 10362
rect 3413 10310 3415 10362
rect 3169 10308 3175 10310
rect 3231 10308 3255 10310
rect 3311 10308 3335 10310
rect 3391 10308 3415 10310
rect 3471 10308 3477 10310
rect 3169 10299 3477 10308
rect 1584 10192 1636 10198
rect 1582 10160 1584 10169
rect 1636 10160 1638 10169
rect 1582 10095 1638 10104
rect 5388 9820 5696 9829
rect 5388 9818 5394 9820
rect 5450 9818 5474 9820
rect 5530 9818 5554 9820
rect 5610 9818 5634 9820
rect 5690 9818 5696 9820
rect 5450 9766 5452 9818
rect 5632 9766 5634 9818
rect 5388 9764 5394 9766
rect 5450 9764 5474 9766
rect 5530 9764 5554 9766
rect 5610 9764 5634 9766
rect 5690 9764 5696 9766
rect 5388 9755 5696 9764
rect 6840 9450 6868 14758
rect 7024 14618 7052 19200
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7576 17241 7604 17274
rect 7562 17232 7618 17241
rect 7380 17196 7432 17202
rect 7562 17167 7618 17176
rect 7380 17138 7432 17144
rect 7392 17105 7420 17138
rect 7378 17096 7434 17105
rect 7760 17082 7788 19200
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 8128 17270 8156 17818
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8116 17264 8168 17270
rect 8300 17264 8352 17270
rect 8116 17206 8168 17212
rect 8298 17232 8300 17241
rect 8352 17232 8354 17241
rect 7760 17054 7972 17082
rect 7378 17031 7434 17040
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 16454 7144 16934
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7116 16238 7328 16266
rect 7116 16182 7144 16238
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 7196 16176 7248 16182
rect 7196 16118 7248 16124
rect 7208 15858 7236 16118
rect 7116 15830 7236 15858
rect 7116 15706 7144 15830
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7104 15496 7156 15502
rect 7208 15484 7236 15642
rect 7156 15456 7236 15484
rect 7104 15438 7156 15444
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7116 13326 7144 15438
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7208 14346 7236 14962
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7300 13870 7328 16238
rect 7392 15638 7420 17031
rect 7608 16892 7916 16901
rect 7608 16890 7614 16892
rect 7670 16890 7694 16892
rect 7750 16890 7774 16892
rect 7830 16890 7854 16892
rect 7910 16890 7916 16892
rect 7670 16838 7672 16890
rect 7852 16838 7854 16890
rect 7608 16836 7614 16838
rect 7670 16836 7694 16838
rect 7750 16836 7774 16838
rect 7830 16836 7854 16838
rect 7910 16836 7916 16838
rect 7608 16827 7916 16836
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7760 16017 7788 16050
rect 7852 16046 7880 16458
rect 7840 16040 7892 16046
rect 7746 16008 7802 16017
rect 7840 15982 7892 15988
rect 7746 15943 7802 15952
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7484 13802 7512 15846
rect 7608 15804 7916 15813
rect 7608 15802 7614 15804
rect 7670 15802 7694 15804
rect 7750 15802 7774 15804
rect 7830 15802 7854 15804
rect 7910 15802 7916 15804
rect 7670 15750 7672 15802
rect 7852 15750 7854 15802
rect 7608 15748 7614 15750
rect 7670 15748 7694 15750
rect 7750 15748 7774 15750
rect 7830 15748 7854 15750
rect 7910 15748 7916 15750
rect 7608 15739 7916 15748
rect 7944 15162 7972 17054
rect 8128 16794 8156 17206
rect 8298 17167 8354 17176
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8404 16794 8432 17070
rect 8496 16998 8524 17546
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8588 17105 8616 17138
rect 8574 17096 8630 17105
rect 8630 17054 8800 17082
rect 9232 17066 9260 19200
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 8574 17031 8630 17040
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 8036 15706 8064 16526
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7930 14920 7986 14929
rect 7930 14855 7986 14864
rect 7608 14716 7916 14725
rect 7608 14714 7614 14716
rect 7670 14714 7694 14716
rect 7750 14714 7774 14716
rect 7830 14714 7854 14716
rect 7910 14714 7916 14716
rect 7670 14662 7672 14714
rect 7852 14662 7854 14714
rect 7608 14660 7614 14662
rect 7670 14660 7694 14662
rect 7750 14660 7774 14662
rect 7830 14660 7854 14662
rect 7910 14660 7916 14662
rect 7608 14651 7916 14660
rect 7944 14618 7972 14855
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7608 13628 7916 13637
rect 7608 13626 7614 13628
rect 7670 13626 7694 13628
rect 7750 13626 7774 13628
rect 7830 13626 7854 13628
rect 7910 13626 7916 13628
rect 7670 13574 7672 13626
rect 7852 13574 7854 13626
rect 7608 13572 7614 13574
rect 7670 13572 7694 13574
rect 7750 13572 7774 13574
rect 7830 13572 7854 13574
rect 7910 13572 7916 13574
rect 7608 13563 7916 13572
rect 7104 13320 7156 13326
rect 8036 13297 8064 15438
rect 8128 15026 8156 16730
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8312 16289 8340 16526
rect 8404 16454 8432 16730
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8298 16280 8354 16289
rect 8298 16215 8354 16224
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8220 14550 8248 15846
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8312 14278 8340 16050
rect 8496 15638 8524 16934
rect 8772 16658 8800 17054
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 7104 13262 7156 13268
rect 8022 13288 8078 13297
rect 8022 13223 8078 13232
rect 8404 13190 8432 14350
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8496 12646 8524 15574
rect 8588 14618 8616 16186
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8668 16040 8720 16046
rect 8666 16008 8668 16017
rect 8944 16040 8996 16046
rect 8720 16008 8722 16017
rect 8666 15943 8722 15952
rect 8942 16008 8944 16017
rect 8996 16008 8998 16017
rect 8942 15943 8998 15952
rect 8680 15638 8708 15943
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 9048 15366 9076 16050
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8758 15056 8814 15065
rect 8864 15026 8892 15302
rect 8758 14991 8814 15000
rect 8852 15020 8904 15026
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8772 13938 8800 14991
rect 8852 14962 8904 14968
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9048 12714 9076 14758
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 7608 12540 7916 12549
rect 7608 12538 7614 12540
rect 7670 12538 7694 12540
rect 7750 12538 7774 12540
rect 7830 12538 7854 12540
rect 7910 12538 7916 12540
rect 7670 12486 7672 12538
rect 7852 12486 7854 12538
rect 7608 12484 7614 12486
rect 7670 12484 7694 12486
rect 7750 12484 7774 12486
rect 7830 12484 7854 12486
rect 7910 12484 7916 12486
rect 7608 12475 7916 12484
rect 9140 11801 9168 16934
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 16153 9352 16390
rect 9310 16144 9366 16153
rect 9310 16079 9366 16088
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9232 13938 9260 15506
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9324 12986 9352 16079
rect 9416 16046 9444 17682
rect 9692 17082 9720 19230
rect 9876 19122 9904 19230
rect 9954 19200 10010 20000
rect 10690 19200 10746 20000
rect 11426 19200 11482 20000
rect 11808 19230 12112 19258
rect 9968 19122 9996 19200
rect 9876 19094 9996 19122
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 9827 17436 10135 17445
rect 9827 17434 9833 17436
rect 9889 17434 9913 17436
rect 9969 17434 9993 17436
rect 10049 17434 10073 17436
rect 10129 17434 10135 17436
rect 9889 17382 9891 17434
rect 10071 17382 10073 17434
rect 9827 17380 9833 17382
rect 9889 17380 9913 17382
rect 9969 17380 9993 17382
rect 10049 17380 10073 17382
rect 10129 17380 10135 17382
rect 9827 17371 10135 17380
rect 9692 17054 9812 17082
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9494 16280 9550 16289
rect 9494 16215 9550 16224
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9416 15502 9444 15982
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9508 14385 9536 16215
rect 9600 14958 9628 16390
rect 9692 15570 9720 16934
rect 9784 16522 9812 17054
rect 10244 16998 10272 17546
rect 10428 17202 10456 17818
rect 11072 17202 11192 17218
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 11060 17196 11192 17202
rect 11112 17190 11192 17196
rect 11060 17138 11112 17144
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10244 16833 10272 16934
rect 10230 16824 10286 16833
rect 10048 16788 10100 16794
rect 10230 16759 10232 16768
rect 10048 16730 10100 16736
rect 10284 16759 10286 16768
rect 10324 16788 10376 16794
rect 10232 16730 10284 16736
rect 10324 16730 10376 16736
rect 10060 16658 10088 16730
rect 10244 16699 10272 16730
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9827 16348 10135 16357
rect 9827 16346 9833 16348
rect 9889 16346 9913 16348
rect 9969 16346 9993 16348
rect 10049 16346 10073 16348
rect 10129 16346 10135 16348
rect 9889 16294 9891 16346
rect 10071 16294 10073 16346
rect 9827 16292 9833 16294
rect 9889 16292 9913 16294
rect 9969 16292 9993 16294
rect 10049 16292 10073 16294
rect 10129 16292 10135 16294
rect 9827 16283 10135 16292
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9772 15632 9824 15638
rect 9770 15600 9772 15609
rect 9824 15600 9826 15609
rect 9680 15564 9732 15570
rect 9770 15535 9826 15544
rect 9680 15506 9732 15512
rect 9968 15473 9996 16118
rect 9954 15464 10010 15473
rect 9954 15399 10010 15408
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9494 14376 9550 14385
rect 9494 14311 9550 14320
rect 9402 13968 9458 13977
rect 9402 13903 9404 13912
rect 9456 13903 9458 13912
rect 9404 13874 9456 13880
rect 9508 13818 9536 14311
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9600 14074 9628 14214
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9692 13938 9720 15302
rect 9827 15260 10135 15269
rect 9827 15258 9833 15260
rect 9889 15258 9913 15260
rect 9969 15258 9993 15260
rect 10049 15258 10073 15260
rect 10129 15258 10135 15260
rect 9889 15206 9891 15258
rect 10071 15206 10073 15258
rect 9827 15204 9833 15206
rect 9889 15204 9913 15206
rect 9969 15204 9993 15206
rect 10049 15204 10073 15206
rect 10129 15204 10135 15206
rect 9827 15195 10135 15204
rect 10336 14958 10364 16730
rect 10428 16590 10456 17138
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10784 16992 10836 16998
rect 10612 16952 10784 16980
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10612 16522 10640 16952
rect 10784 16934 10836 16940
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10506 16280 10562 16289
rect 10506 16215 10562 16224
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15026 10456 15846
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14346 10088 14758
rect 10138 14648 10194 14657
rect 10138 14583 10194 14592
rect 10152 14550 10180 14583
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 9827 14172 10135 14181
rect 9827 14170 9833 14172
rect 9889 14170 9913 14172
rect 9969 14170 9993 14172
rect 10049 14170 10073 14172
rect 10129 14170 10135 14172
rect 9889 14118 9891 14170
rect 10071 14118 10073 14170
rect 9827 14116 9833 14118
rect 9889 14116 9913 14118
rect 9969 14116 9993 14118
rect 10049 14116 10073 14118
rect 10129 14116 10135 14118
rect 9827 14107 10135 14116
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10060 13841 10088 13874
rect 10046 13832 10102 13841
rect 9508 13790 9904 13818
rect 9876 13326 9904 13790
rect 10046 13767 10102 13776
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9827 13084 10135 13093
rect 9827 13082 9833 13084
rect 9889 13082 9913 13084
rect 9969 13082 9993 13084
rect 10049 13082 10073 13084
rect 10129 13082 10135 13084
rect 9889 13030 9891 13082
rect 10071 13030 10073 13082
rect 9827 13028 9833 13030
rect 9889 13028 9913 13030
rect 9969 13028 9993 13030
rect 10049 13028 10073 13030
rect 10129 13028 10135 13030
rect 9827 13019 10135 13028
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9827 11996 10135 12005
rect 9827 11994 9833 11996
rect 9889 11994 9913 11996
rect 9969 11994 9993 11996
rect 10049 11994 10073 11996
rect 10129 11994 10135 11996
rect 9889 11942 9891 11994
rect 10071 11942 10073 11994
rect 9827 11940 9833 11942
rect 9889 11940 9913 11942
rect 9969 11940 9993 11942
rect 10049 11940 10073 11942
rect 10129 11940 10135 11942
rect 9827 11931 10135 11940
rect 9126 11792 9182 11801
rect 9126 11727 9182 11736
rect 10244 11694 10272 14826
rect 10324 14612 10376 14618
rect 10376 14572 10456 14600
rect 10324 14554 10376 14560
rect 10322 14512 10378 14521
rect 10322 14447 10378 14456
rect 10336 13870 10364 14447
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10324 13728 10376 13734
rect 10428 13716 10456 14572
rect 10520 14006 10548 16215
rect 10612 15201 10640 16458
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10598 15192 10654 15201
rect 10598 15127 10654 15136
rect 10612 15026 10640 15127
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10612 13938 10640 14418
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10376 13688 10456 13716
rect 10508 13728 10560 13734
rect 10506 13696 10508 13705
rect 10560 13696 10562 13705
rect 10324 13670 10376 13676
rect 10336 11830 10364 13670
rect 10506 13631 10562 13640
rect 10414 13560 10470 13569
rect 10414 13495 10470 13504
rect 10428 13190 10456 13495
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10520 13025 10548 13398
rect 10612 13326 10640 13874
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10506 13016 10562 13025
rect 10506 12951 10562 12960
rect 10506 12880 10562 12889
rect 10506 12815 10508 12824
rect 10560 12815 10562 12824
rect 10508 12786 10560 12792
rect 10612 12730 10640 13262
rect 10704 12753 10732 16390
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10796 15570 10824 16050
rect 10888 15910 10916 16934
rect 10966 16824 11022 16833
rect 10966 16759 11022 16768
rect 10980 16590 11008 16759
rect 11072 16697 11100 17002
rect 11058 16688 11114 16697
rect 11058 16623 11060 16632
rect 11112 16623 11114 16632
rect 11060 16594 11112 16600
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10796 14822 10824 14962
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10874 14648 10930 14657
rect 10874 14583 10930 14592
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 13705 10824 14350
rect 10888 13938 10916 14583
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10782 13696 10838 13705
rect 10782 13631 10838 13640
rect 10428 12702 10640 12730
rect 10690 12744 10746 12753
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 7608 11452 7916 11461
rect 7608 11450 7614 11452
rect 7670 11450 7694 11452
rect 7750 11450 7774 11452
rect 7830 11450 7854 11452
rect 7910 11450 7916 11452
rect 7670 11398 7672 11450
rect 7852 11398 7854 11450
rect 7608 11396 7614 11398
rect 7670 11396 7694 11398
rect 7750 11396 7774 11398
rect 7830 11396 7854 11398
rect 7910 11396 7916 11398
rect 7608 11387 7916 11396
rect 10428 11218 10456 12702
rect 10690 12679 10746 12688
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10520 12374 10548 12582
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10796 11626 10824 13631
rect 10888 11898 10916 13874
rect 10980 12714 11008 16050
rect 11164 15638 11192 17190
rect 11440 16946 11468 19200
rect 11808 17338 11836 19230
rect 12084 19122 12112 19230
rect 12162 19200 12218 20000
rect 12898 19200 12954 20000
rect 13634 19200 13690 20000
rect 14370 19200 14426 20000
rect 15106 19200 15162 20000
rect 15842 19200 15898 20000
rect 16578 19200 16634 20000
rect 16684 19230 16988 19258
rect 12176 19122 12204 19200
rect 12084 19094 12204 19122
rect 13648 17542 13676 19200
rect 14384 18034 14412 19200
rect 15658 19000 15714 19009
rect 15658 18935 15714 18944
rect 14200 18006 14412 18034
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 12992 17264 13044 17270
rect 12992 17206 13044 17212
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 11256 16918 11468 16946
rect 11256 15706 11284 16918
rect 12047 16892 12355 16901
rect 12047 16890 12053 16892
rect 12109 16890 12133 16892
rect 12189 16890 12213 16892
rect 12269 16890 12293 16892
rect 12349 16890 12355 16892
rect 12109 16838 12111 16890
rect 12291 16838 12293 16890
rect 12047 16836 12053 16838
rect 12109 16836 12133 16838
rect 12189 16836 12213 16838
rect 12269 16836 12293 16838
rect 12349 16836 12355 16838
rect 12047 16827 12355 16836
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11152 15632 11204 15638
rect 11204 15580 11284 15586
rect 11152 15574 11284 15580
rect 11164 15558 11284 15574
rect 11058 15328 11114 15337
rect 11058 15263 11114 15272
rect 11072 15026 11100 15263
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11072 14414 11100 14962
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11058 14240 11114 14249
rect 11058 14175 11114 14184
rect 11072 13530 11100 14175
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11164 13326 11192 14758
rect 11256 14346 11284 15558
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11242 14104 11298 14113
rect 11242 14039 11298 14048
rect 11256 14006 11284 14039
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11244 13864 11296 13870
rect 11242 13832 11244 13841
rect 11296 13832 11298 13841
rect 11242 13767 11298 13776
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 13462 11284 13670
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11152 12980 11204 12986
rect 11256 12968 11284 13262
rect 11204 12940 11284 12968
rect 11152 12922 11204 12928
rect 11058 12880 11114 12889
rect 11058 12815 11060 12824
rect 11112 12815 11114 12824
rect 11060 12786 11112 12792
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 11256 12102 11284 12940
rect 11348 12442 11376 16526
rect 11888 16448 11940 16454
rect 11426 16416 11482 16425
rect 12268 16425 12296 16594
rect 11888 16390 11940 16396
rect 12254 16416 12310 16425
rect 11426 16351 11482 16360
rect 11440 14550 11468 16351
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11808 15638 11836 16050
rect 11900 16046 11928 16390
rect 12254 16351 12310 16360
rect 12360 16289 12388 16594
rect 12346 16280 12402 16289
rect 12346 16215 12402 16224
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 11532 14618 11560 14826
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11336 12436 11388 12442
rect 11440 12434 11468 14282
rect 11532 12714 11560 14418
rect 11624 13841 11652 15098
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 14618 11744 14894
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11808 14482 11836 15574
rect 11900 14958 11928 15982
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12047 15804 12355 15813
rect 12047 15802 12053 15804
rect 12109 15802 12133 15804
rect 12189 15802 12213 15804
rect 12269 15802 12293 15804
rect 12349 15802 12355 15804
rect 12109 15750 12111 15802
rect 12291 15750 12293 15802
rect 12047 15748 12053 15750
rect 12109 15748 12133 15750
rect 12189 15748 12213 15750
rect 12269 15748 12293 15750
rect 12349 15748 12355 15750
rect 12047 15739 12355 15748
rect 12452 15706 12480 15846
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12544 15162 12572 15846
rect 12714 15464 12770 15473
rect 12714 15399 12770 15408
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 15162 12664 15302
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11610 13832 11666 13841
rect 11610 13767 11666 13776
rect 11610 13560 11666 13569
rect 11610 13495 11666 13504
rect 11624 13462 11652 13495
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12730 11652 13262
rect 11716 12850 11744 14214
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11520 12708 11572 12714
rect 11624 12702 11744 12730
rect 11520 12650 11572 12656
rect 11440 12406 11652 12434
rect 11336 12378 11388 12384
rect 11624 12306 11652 12406
rect 11716 12345 11744 12702
rect 11702 12336 11758 12345
rect 11612 12300 11664 12306
rect 11702 12271 11758 12280
rect 11612 12242 11664 12248
rect 11808 12238 11836 13670
rect 11900 13326 11928 14894
rect 12047 14716 12355 14725
rect 12047 14714 12053 14716
rect 12109 14714 12133 14716
rect 12189 14714 12213 14716
rect 12269 14714 12293 14716
rect 12349 14714 12355 14716
rect 12109 14662 12111 14714
rect 12291 14662 12293 14714
rect 12047 14660 12053 14662
rect 12109 14660 12133 14662
rect 12189 14660 12213 14662
rect 12269 14660 12293 14662
rect 12349 14660 12355 14662
rect 12047 14651 12355 14660
rect 12254 14512 12310 14521
rect 12254 14447 12310 14456
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 14006 12020 14214
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 12268 13938 12296 14447
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12346 13832 12402 13841
rect 12452 13818 12480 15030
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12530 13832 12586 13841
rect 12452 13790 12530 13818
rect 12346 13767 12402 13776
rect 12530 13767 12586 13776
rect 12360 13716 12388 13767
rect 12360 13688 12480 13716
rect 12047 13628 12355 13637
rect 12047 13626 12053 13628
rect 12109 13626 12133 13628
rect 12189 13626 12213 13628
rect 12269 13626 12293 13628
rect 12349 13626 12355 13628
rect 12109 13574 12111 13626
rect 12291 13574 12293 13626
rect 12047 13572 12053 13574
rect 12109 13572 12133 13574
rect 12189 13572 12213 13574
rect 12269 13572 12293 13574
rect 12349 13572 12355 13574
rect 12047 13563 12355 13572
rect 12164 13524 12216 13530
rect 12452 13512 12480 13688
rect 12636 13569 12664 14010
rect 12164 13466 12216 13472
rect 12360 13484 12480 13512
rect 12622 13560 12678 13569
rect 12622 13495 12678 13504
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11992 13190 12020 13398
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11900 12918 11928 13126
rect 11888 12912 11940 12918
rect 12176 12889 12204 13466
rect 12360 13258 12388 13484
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 11888 12854 11940 12860
rect 12162 12880 12218 12889
rect 12452 12850 12480 13126
rect 12544 12850 12572 13398
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12162 12815 12218 12824
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12636 12714 12664 13262
rect 12728 12986 12756 15399
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12820 12782 12848 17070
rect 13004 15570 13032 17206
rect 13740 17202 13768 17682
rect 14200 17338 14228 18006
rect 14648 17808 14700 17814
rect 14648 17750 14700 17756
rect 14266 17436 14574 17445
rect 14266 17434 14272 17436
rect 14328 17434 14352 17436
rect 14408 17434 14432 17436
rect 14488 17434 14512 17436
rect 14568 17434 14574 17436
rect 14328 17382 14330 17434
rect 14510 17382 14512 17434
rect 14266 17380 14272 17382
rect 14328 17380 14352 17382
rect 14408 17380 14432 17382
rect 14488 17380 14512 17382
rect 14568 17380 14574 17382
rect 14266 17371 14574 17380
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13740 17082 13768 17138
rect 14188 17128 14240 17134
rect 13464 16794 13492 17070
rect 13740 17054 13952 17082
rect 14188 17070 14240 17076
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13634 16688 13690 16697
rect 13634 16623 13690 16632
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13556 16454 13584 16526
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13188 16114 13216 16390
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13188 15745 13216 16050
rect 13174 15736 13230 15745
rect 13174 15671 13230 15680
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12912 14074 12940 15098
rect 13004 14958 13032 15506
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13004 14346 13032 14894
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14521 13124 14758
rect 13082 14512 13138 14521
rect 13082 14447 13138 14456
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13084 14272 13136 14278
rect 13082 14240 13084 14249
rect 13136 14240 13138 14249
rect 13082 14175 13138 14184
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12912 13841 12940 13874
rect 12898 13832 12954 13841
rect 12898 13767 12954 13776
rect 12898 13696 12954 13705
rect 12898 13631 12954 13640
rect 12912 13190 12940 13631
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 11900 11354 11928 12582
rect 12047 12540 12355 12549
rect 12047 12538 12053 12540
rect 12109 12538 12133 12540
rect 12189 12538 12213 12540
rect 12269 12538 12293 12540
rect 12349 12538 12355 12540
rect 12109 12486 12111 12538
rect 12291 12486 12293 12538
rect 12047 12484 12053 12486
rect 12109 12484 12133 12486
rect 12189 12484 12213 12486
rect 12269 12484 12293 12486
rect 12349 12484 12355 12486
rect 12047 12475 12355 12484
rect 12622 12472 12678 12481
rect 12622 12407 12678 12416
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 11558 12296 12174
rect 12636 11762 12664 12407
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12256 11552 12308 11558
rect 13004 11529 13032 13942
rect 13096 13274 13124 14010
rect 13188 13394 13216 15370
rect 13280 14793 13308 16186
rect 13358 15872 13414 15881
rect 13358 15807 13414 15816
rect 13266 14784 13322 14793
rect 13266 14719 13322 14728
rect 13266 14512 13322 14521
rect 13266 14447 13322 14456
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13096 13246 13216 13274
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13096 12306 13124 12786
rect 13188 12434 13216 13246
rect 13280 13138 13308 14447
rect 13372 13734 13400 15807
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13358 13424 13414 13433
rect 13464 13394 13492 14418
rect 13556 14006 13584 15098
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13358 13359 13360 13368
rect 13412 13359 13414 13368
rect 13452 13388 13504 13394
rect 13360 13330 13412 13336
rect 13452 13330 13504 13336
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13280 13110 13400 13138
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13280 12782 13308 12922
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13372 12481 13400 13110
rect 13358 12472 13414 12481
rect 13188 12406 13308 12434
rect 13358 12407 13414 12416
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13280 12238 13308 12406
rect 13452 12368 13504 12374
rect 13358 12336 13414 12345
rect 13452 12310 13504 12316
rect 13358 12271 13414 12280
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13372 11778 13400 12271
rect 13280 11762 13400 11778
rect 13268 11756 13400 11762
rect 13320 11750 13400 11756
rect 13268 11698 13320 11704
rect 13464 11665 13492 12310
rect 13450 11656 13506 11665
rect 13450 11591 13506 11600
rect 12256 11494 12308 11500
rect 12990 11520 13046 11529
rect 12047 11452 12355 11461
rect 12990 11455 13046 11464
rect 12047 11450 12053 11452
rect 12109 11450 12133 11452
rect 12189 11450 12213 11452
rect 12269 11450 12293 11452
rect 12349 11450 12355 11452
rect 12109 11398 12111 11450
rect 12291 11398 12293 11450
rect 12047 11396 12053 11398
rect 12109 11396 12133 11398
rect 12189 11396 12213 11398
rect 12269 11396 12293 11398
rect 12349 11396 12355 11398
rect 12047 11387 12355 11396
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 13556 11098 13584 13262
rect 13464 11082 13584 11098
rect 13452 11076 13584 11082
rect 13504 11070 13584 11076
rect 13452 11018 13504 11024
rect 9827 10908 10135 10917
rect 9827 10906 9833 10908
rect 9889 10906 9913 10908
rect 9969 10906 9993 10908
rect 10049 10906 10073 10908
rect 10129 10906 10135 10908
rect 9889 10854 9891 10906
rect 10071 10854 10073 10906
rect 9827 10852 9833 10854
rect 9889 10852 9913 10854
rect 9969 10852 9993 10854
rect 10049 10852 10073 10854
rect 10129 10852 10135 10854
rect 9827 10843 10135 10852
rect 7608 10364 7916 10373
rect 7608 10362 7614 10364
rect 7670 10362 7694 10364
rect 7750 10362 7774 10364
rect 7830 10362 7854 10364
rect 7910 10362 7916 10364
rect 7670 10310 7672 10362
rect 7852 10310 7854 10362
rect 7608 10308 7614 10310
rect 7670 10308 7694 10310
rect 7750 10308 7774 10310
rect 7830 10308 7854 10310
rect 7910 10308 7916 10310
rect 7608 10299 7916 10308
rect 12047 10364 12355 10373
rect 12047 10362 12053 10364
rect 12109 10362 12133 10364
rect 12189 10362 12213 10364
rect 12269 10362 12293 10364
rect 12349 10362 12355 10364
rect 12109 10310 12111 10362
rect 12291 10310 12293 10362
rect 12047 10308 12053 10310
rect 12109 10308 12133 10310
rect 12189 10308 12213 10310
rect 12269 10308 12293 10310
rect 12349 10308 12355 10310
rect 12047 10299 12355 10308
rect 13648 10062 13676 16623
rect 13740 13462 13768 16934
rect 13924 16794 13952 17054
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16250 13860 16390
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13818 15736 13874 15745
rect 13818 15671 13874 15680
rect 13832 15502 13860 15671
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13832 15162 13860 15438
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13924 14482 13952 16730
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 14016 15366 14044 16458
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 14002 15192 14058 15201
rect 14200 15178 14228 17070
rect 14292 16590 14320 17274
rect 14660 17241 14688 17750
rect 14740 17264 14792 17270
rect 14646 17232 14702 17241
rect 14740 17206 14792 17212
rect 14646 17167 14702 17176
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14266 16348 14574 16357
rect 14266 16346 14272 16348
rect 14328 16346 14352 16348
rect 14408 16346 14432 16348
rect 14488 16346 14512 16348
rect 14568 16346 14574 16348
rect 14328 16294 14330 16346
rect 14510 16294 14512 16346
rect 14266 16292 14272 16294
rect 14328 16292 14352 16294
rect 14408 16292 14432 16294
rect 14488 16292 14512 16294
rect 14568 16292 14574 16294
rect 14266 16283 14574 16292
rect 14660 16096 14688 16934
rect 14752 16454 14780 17206
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14740 16448 14792 16454
rect 14936 16402 14964 16594
rect 14740 16390 14792 16396
rect 14752 16114 14780 16390
rect 14844 16374 14964 16402
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 14568 16068 14688 16096
rect 14740 16108 14792 16114
rect 14568 15570 14596 16068
rect 14740 16050 14792 16056
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14266 15260 14574 15269
rect 14266 15258 14272 15260
rect 14328 15258 14352 15260
rect 14408 15258 14432 15260
rect 14488 15258 14512 15260
rect 14568 15258 14574 15260
rect 14328 15206 14330 15258
rect 14510 15206 14512 15258
rect 14266 15204 14272 15206
rect 14328 15204 14352 15206
rect 14408 15204 14432 15206
rect 14488 15204 14512 15206
rect 14568 15204 14574 15206
rect 14266 15195 14574 15204
rect 14002 15127 14058 15136
rect 14108 15150 14228 15178
rect 13912 14476 13964 14482
rect 13832 14436 13912 14464
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13832 13326 13860 14436
rect 13912 14418 13964 14424
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 12776 13780 12782
rect 13832 12764 13860 13262
rect 13780 12736 13860 12764
rect 13728 12718 13780 12724
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 12442 13860 12582
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13726 12336 13782 12345
rect 13726 12271 13782 12280
rect 13820 12300 13872 12306
rect 13740 11150 13768 12271
rect 13820 12242 13872 12248
rect 13832 12102 13860 12242
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13818 11928 13874 11937
rect 13924 11898 13952 14282
rect 14016 13870 14044 15127
rect 14108 14906 14136 15150
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14108 14878 14228 14906
rect 14094 14784 14150 14793
rect 14094 14719 14150 14728
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14002 13560 14058 13569
rect 14002 13495 14058 13504
rect 14016 12209 14044 13495
rect 14108 12442 14136 14719
rect 14200 12986 14228 14878
rect 14384 14793 14412 15030
rect 14370 14784 14426 14793
rect 14370 14719 14426 14728
rect 14660 14482 14688 15914
rect 14752 14793 14780 16050
rect 14844 16046 14872 16374
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14738 14784 14794 14793
rect 14738 14719 14794 14728
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14266 14172 14574 14181
rect 14266 14170 14272 14172
rect 14328 14170 14352 14172
rect 14408 14170 14432 14172
rect 14488 14170 14512 14172
rect 14568 14170 14574 14172
rect 14328 14118 14330 14170
rect 14510 14118 14512 14170
rect 14266 14116 14272 14118
rect 14328 14116 14352 14118
rect 14408 14116 14432 14118
rect 14488 14116 14512 14118
rect 14568 14116 14574 14118
rect 14266 14107 14574 14116
rect 14648 13864 14700 13870
rect 14700 13812 14780 13818
rect 14648 13806 14780 13812
rect 14660 13790 14780 13806
rect 14266 13084 14574 13093
rect 14266 13082 14272 13084
rect 14328 13082 14352 13084
rect 14408 13082 14432 13084
rect 14488 13082 14512 13084
rect 14568 13082 14574 13084
rect 14328 13030 14330 13082
rect 14510 13030 14512 13082
rect 14266 13028 14272 13030
rect 14328 13028 14352 13030
rect 14408 13028 14432 13030
rect 14488 13028 14512 13030
rect 14568 13028 14574 13030
rect 14266 13019 14574 13028
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14646 12880 14702 12889
rect 14646 12815 14702 12824
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14188 12232 14240 12238
rect 14002 12200 14058 12209
rect 14188 12174 14240 12180
rect 14002 12135 14058 12144
rect 13818 11863 13874 11872
rect 13912 11892 13964 11898
rect 13832 11694 13860 11863
rect 13912 11834 13964 11840
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 14016 10674 14044 12135
rect 14200 10810 14228 12174
rect 14266 11996 14574 12005
rect 14266 11994 14272 11996
rect 14328 11994 14352 11996
rect 14408 11994 14432 11996
rect 14488 11994 14512 11996
rect 14568 11994 14574 11996
rect 14328 11942 14330 11994
rect 14510 11942 14512 11994
rect 14266 11940 14272 11942
rect 14328 11940 14352 11942
rect 14408 11940 14432 11942
rect 14488 11940 14512 11942
rect 14568 11940 14574 11942
rect 14266 11931 14574 11940
rect 14660 11830 14688 12815
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14476 11529 14504 11698
rect 14462 11520 14518 11529
rect 14462 11455 14518 11464
rect 14278 11384 14334 11393
rect 14278 11319 14280 11328
rect 14332 11319 14334 11328
rect 14280 11290 14332 11296
rect 14660 11218 14688 11766
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14266 10908 14574 10917
rect 14266 10906 14272 10908
rect 14328 10906 14352 10908
rect 14408 10906 14432 10908
rect 14488 10906 14512 10908
rect 14568 10906 14574 10908
rect 14328 10854 14330 10906
rect 14510 10854 14512 10906
rect 14266 10852 14272 10854
rect 14328 10852 14352 10854
rect 14408 10852 14432 10854
rect 14488 10852 14512 10854
rect 14568 10852 14574 10854
rect 14266 10843 14574 10852
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14752 10130 14780 13790
rect 14844 13433 14872 15438
rect 14936 15094 14964 16118
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15028 15609 15056 15982
rect 15014 15600 15070 15609
rect 15014 15535 15016 15544
rect 15068 15535 15070 15544
rect 15198 15600 15254 15609
rect 15198 15535 15254 15544
rect 15016 15506 15068 15512
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15028 15337 15056 15370
rect 15014 15328 15070 15337
rect 15014 15263 15070 15272
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 14922 14784 14978 14793
rect 14922 14719 14978 14728
rect 14936 14113 14964 14719
rect 15028 14482 15056 14962
rect 15212 14521 15240 15535
rect 15290 15328 15346 15337
rect 15290 15263 15346 15272
rect 15304 14890 15332 15263
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15198 14512 15254 14521
rect 15016 14476 15068 14482
rect 15198 14447 15254 14456
rect 15016 14418 15068 14424
rect 15106 14376 15162 14385
rect 15304 14346 15332 14826
rect 15106 14311 15162 14320
rect 15292 14340 15344 14346
rect 14922 14104 14978 14113
rect 15120 14074 15148 14311
rect 15292 14282 15344 14288
rect 14922 14039 14978 14048
rect 15108 14068 15160 14074
rect 14936 14006 14964 14039
rect 15108 14010 15160 14016
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15108 13728 15160 13734
rect 15212 13705 15240 13942
rect 15108 13670 15160 13676
rect 15198 13696 15254 13705
rect 14830 13424 14886 13433
rect 14830 13359 14886 13368
rect 14844 12306 14872 13359
rect 15014 13152 15070 13161
rect 15014 13087 15070 13096
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14936 12306 14964 12922
rect 15028 12442 15056 13087
rect 15120 12889 15148 13670
rect 15198 13631 15254 13640
rect 15106 12880 15162 12889
rect 15106 12815 15162 12824
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14830 12200 14886 12209
rect 14830 12135 14886 12144
rect 14924 12164 14976 12170
rect 14844 10742 14872 12135
rect 14924 12106 14976 12112
rect 14936 12073 14964 12106
rect 14922 12064 14978 12073
rect 14922 11999 14978 12008
rect 15028 11218 15056 12378
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 15028 10470 15056 11154
rect 15120 10810 15148 12242
rect 15212 11762 15240 13631
rect 15304 13258 15332 14282
rect 15396 13802 15424 15982
rect 15488 15162 15516 16390
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15488 14657 15516 15098
rect 15474 14648 15530 14657
rect 15474 14583 15530 14592
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 15292 13252 15344 13258
rect 15344 13212 15424 13240
rect 15292 13194 15344 13200
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15304 12714 15332 12854
rect 15396 12850 15424 13212
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15396 12594 15424 12786
rect 15304 12566 15424 12594
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15304 11354 15332 12566
rect 15488 12458 15516 14583
rect 15580 13938 15608 15642
rect 15672 14929 15700 18935
rect 15856 17898 15884 19200
rect 16592 19122 16620 19200
rect 16684 19122 16712 19230
rect 16592 19094 16712 19122
rect 15856 17870 15976 17898
rect 15842 16280 15898 16289
rect 15842 16215 15844 16224
rect 15896 16215 15898 16224
rect 15844 16186 15896 16192
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15752 15496 15804 15502
rect 15856 15473 15884 16050
rect 15752 15438 15804 15444
rect 15842 15464 15898 15473
rect 15658 14920 15714 14929
rect 15658 14855 15714 14864
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15672 13870 15700 14554
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12646 15608 12786
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15396 12430 15516 12458
rect 15396 11558 15424 12430
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15488 12084 15516 12310
rect 15580 12238 15608 12582
rect 15672 12442 15700 13806
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15568 12232 15620 12238
rect 15566 12200 15568 12209
rect 15660 12232 15712 12238
rect 15620 12200 15622 12209
rect 15764 12220 15792 15438
rect 15842 15399 15898 15408
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15856 13841 15884 13874
rect 15842 13832 15898 13841
rect 15842 13767 15898 13776
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15712 12192 15792 12220
rect 15660 12174 15712 12180
rect 15566 12135 15622 12144
rect 15488 12056 15700 12084
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15672 11132 15700 12056
rect 15750 12064 15806 12073
rect 15750 11999 15806 12008
rect 15764 11558 15792 11999
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11286 15792 11494
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15752 11144 15804 11150
rect 15672 11112 15752 11132
rect 15804 11112 15806 11121
rect 15672 11104 15750 11112
rect 15750 11047 15806 11056
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15764 10606 15792 11047
rect 15856 10674 15884 13262
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15948 10266 15976 17870
rect 16026 17776 16082 17785
rect 16026 17711 16082 17720
rect 16040 15065 16068 17711
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16132 16590 16160 16730
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16132 15502 16160 16526
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16026 15056 16082 15065
rect 16026 14991 16082 15000
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16040 13530 16068 13942
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 16040 10674 16068 12718
rect 16132 12628 16160 14894
rect 16224 14346 16252 15982
rect 16316 15881 16344 15982
rect 16408 15978 16436 17070
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16486 16892 16794 16901
rect 16486 16890 16492 16892
rect 16548 16890 16572 16892
rect 16628 16890 16652 16892
rect 16708 16890 16732 16892
rect 16788 16890 16794 16892
rect 16548 16838 16550 16890
rect 16730 16838 16732 16890
rect 16486 16836 16492 16838
rect 16548 16836 16572 16838
rect 16628 16836 16652 16838
rect 16708 16836 16732 16838
rect 16788 16836 16794 16838
rect 16486 16827 16794 16836
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16776 16017 16804 16594
rect 16868 16561 16896 16934
rect 16854 16552 16910 16561
rect 16854 16487 16910 16496
rect 16762 16008 16818 16017
rect 16396 15972 16448 15978
rect 16762 15943 16818 15952
rect 16396 15914 16448 15920
rect 16302 15872 16358 15881
rect 16302 15807 16358 15816
rect 16408 14890 16436 15914
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16486 15804 16794 15813
rect 16486 15802 16492 15804
rect 16548 15802 16572 15804
rect 16628 15802 16652 15804
rect 16708 15802 16732 15804
rect 16788 15802 16794 15804
rect 16548 15750 16550 15802
rect 16730 15750 16732 15802
rect 16486 15748 16492 15750
rect 16548 15748 16572 15750
rect 16628 15748 16652 15750
rect 16708 15748 16732 15750
rect 16788 15748 16794 15750
rect 16486 15739 16794 15748
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16224 13870 16252 14282
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16408 13394 16436 14826
rect 16486 14716 16794 14725
rect 16486 14714 16492 14716
rect 16548 14714 16572 14716
rect 16628 14714 16652 14716
rect 16708 14714 16732 14716
rect 16788 14714 16794 14716
rect 16548 14662 16550 14714
rect 16730 14662 16732 14714
rect 16486 14660 16492 14662
rect 16548 14660 16572 14662
rect 16628 14660 16652 14662
rect 16708 14660 16732 14662
rect 16788 14660 16794 14662
rect 16486 14651 16794 14660
rect 16868 14521 16896 15846
rect 16854 14512 16910 14521
rect 16854 14447 16910 14456
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16486 13628 16794 13637
rect 16486 13626 16492 13628
rect 16548 13626 16572 13628
rect 16628 13626 16652 13628
rect 16708 13626 16732 13628
rect 16788 13626 16794 13628
rect 16548 13574 16550 13626
rect 16730 13574 16732 13626
rect 16486 13572 16492 13574
rect 16548 13572 16572 13574
rect 16628 13572 16652 13574
rect 16708 13572 16732 13574
rect 16788 13572 16794 13574
rect 16486 13563 16794 13572
rect 16670 13424 16726 13433
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16396 13388 16448 13394
rect 16670 13359 16726 13368
rect 16396 13330 16448 13336
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16224 12730 16252 13194
rect 16316 12918 16344 13330
rect 16684 13326 16712 13359
rect 16672 13320 16724 13326
rect 16486 13288 16542 13297
rect 16396 13252 16448 13258
rect 16672 13262 16724 13268
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16486 13223 16542 13232
rect 16396 13194 16448 13200
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16408 12850 16436 13194
rect 16500 13190 16528 13223
rect 16488 13184 16540 13190
rect 16776 13161 16804 13262
rect 16488 13126 16540 13132
rect 16762 13152 16818 13161
rect 16762 13087 16818 13096
rect 16486 12880 16542 12889
rect 16396 12844 16448 12850
rect 16486 12815 16542 12824
rect 16396 12786 16448 12792
rect 16224 12714 16344 12730
rect 16224 12708 16356 12714
rect 16224 12702 16304 12708
rect 16304 12650 16356 12656
rect 16132 12600 16252 12628
rect 16118 12472 16174 12481
rect 16118 12407 16174 12416
rect 16132 12306 16160 12407
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16132 11801 16160 12106
rect 16118 11792 16174 11801
rect 16118 11727 16174 11736
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11014 16160 11494
rect 16224 11014 16252 12600
rect 16316 12238 16344 12650
rect 16500 12646 16528 12815
rect 16580 12776 16632 12782
rect 16578 12744 16580 12753
rect 16632 12744 16634 12753
rect 16578 12679 16634 12688
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16486 12540 16794 12549
rect 16486 12538 16492 12540
rect 16548 12538 16572 12540
rect 16628 12538 16652 12540
rect 16708 12538 16732 12540
rect 16788 12538 16794 12540
rect 16548 12486 16550 12538
rect 16730 12486 16732 12538
rect 16486 12484 16492 12486
rect 16548 12484 16572 12486
rect 16628 12484 16652 12486
rect 16708 12484 16732 12486
rect 16788 12484 16794 12486
rect 16486 12475 16794 12484
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11529 16344 12038
rect 16408 11898 16436 12310
rect 16396 11892 16448 11898
rect 16868 11880 16896 14282
rect 16396 11834 16448 11840
rect 16776 11852 16896 11880
rect 16776 11665 16804 11852
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16762 11656 16818 11665
rect 16762 11591 16818 11600
rect 16302 11520 16358 11529
rect 16302 11455 16358 11464
rect 16486 11452 16794 11461
rect 16486 11450 16492 11452
rect 16548 11450 16572 11452
rect 16628 11450 16652 11452
rect 16708 11450 16732 11452
rect 16788 11450 16794 11452
rect 16548 11398 16550 11450
rect 16730 11398 16732 11450
rect 16486 11396 16492 11398
rect 16548 11396 16572 11398
rect 16628 11396 16652 11398
rect 16708 11396 16732 11398
rect 16788 11396 16794 11398
rect 16486 11387 16794 11396
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16408 10198 16436 11086
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10742 16528 11018
rect 16868 10810 16896 11698
rect 16960 11354 16988 19230
rect 17314 19200 17370 20000
rect 18050 19200 18106 20000
rect 18786 19200 18842 20000
rect 18892 19230 19288 19258
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 17052 16182 17080 17206
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17052 14958 17080 16118
rect 17144 14958 17172 17818
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17236 16046 17264 17206
rect 17592 17060 17644 17066
rect 17592 17002 17644 17008
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17236 15094 17264 15982
rect 17328 15434 17356 16458
rect 17604 16182 17632 17002
rect 17592 16176 17644 16182
rect 17592 16118 17644 16124
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17328 15337 17356 15370
rect 17314 15328 17370 15337
rect 17314 15263 17370 15272
rect 17604 15178 17632 16118
rect 18064 15858 18092 19200
rect 18800 19122 18828 19200
rect 18892 19122 18920 19230
rect 18800 19094 18920 19122
rect 18705 17436 19013 17445
rect 18705 17434 18711 17436
rect 18767 17434 18791 17436
rect 18847 17434 18871 17436
rect 18927 17434 18951 17436
rect 19007 17434 19013 17436
rect 18767 17382 18769 17434
rect 18949 17382 18951 17434
rect 18705 17380 18711 17382
rect 18767 17380 18791 17382
rect 18847 17380 18871 17382
rect 18927 17380 18951 17382
rect 19007 17380 19013 17382
rect 18705 17371 19013 17380
rect 19154 17368 19210 17377
rect 19154 17303 19210 17312
rect 19062 17232 19118 17241
rect 18328 17196 18380 17202
rect 19168 17218 19196 17303
rect 19118 17190 19196 17218
rect 19062 17167 19118 17176
rect 18328 17138 18380 17144
rect 18340 16522 18368 17138
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18064 15830 18184 15858
rect 17604 15150 17724 15178
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13530 17080 13670
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17052 13297 17080 13466
rect 17038 13288 17094 13297
rect 17144 13258 17172 13806
rect 17236 13433 17264 13874
rect 17222 13424 17278 13433
rect 17328 13394 17356 13874
rect 17222 13359 17278 13368
rect 17316 13388 17368 13394
rect 17038 13223 17094 13232
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17040 13184 17092 13190
rect 17236 13138 17264 13359
rect 17316 13330 17368 13336
rect 17314 13288 17370 13297
rect 17314 13223 17370 13232
rect 17040 13126 17092 13132
rect 17052 12850 17080 13126
rect 17144 13110 17264 13138
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 17144 11218 17172 13110
rect 17222 13016 17278 13025
rect 17222 12951 17278 12960
rect 17236 12646 17264 12951
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 17144 10742 17172 11154
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17236 10470 17264 12582
rect 17328 12434 17356 13223
rect 17420 12986 17448 14418
rect 17512 13530 17540 14894
rect 17696 14822 17724 15150
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17696 14278 17724 14758
rect 17788 14482 17816 14962
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17512 12866 17540 13330
rect 17696 13258 17724 14214
rect 17788 14113 17816 14282
rect 17774 14104 17830 14113
rect 17774 14039 17830 14048
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17696 13025 17724 13194
rect 17682 13016 17738 13025
rect 17682 12951 17738 12960
rect 17788 12900 17816 14039
rect 17880 14006 17908 15098
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17972 14482 18000 15030
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17972 13852 18000 14418
rect 18064 13977 18092 14758
rect 18050 13968 18106 13977
rect 18050 13903 18106 13912
rect 17880 13824 18000 13852
rect 18050 13832 18106 13841
rect 17880 13530 17908 13824
rect 18050 13767 18106 13776
rect 18064 13734 18092 13767
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17880 13190 17908 13466
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17420 12850 17540 12866
rect 17408 12844 17540 12850
rect 17460 12838 17540 12844
rect 17604 12872 17816 12900
rect 17408 12786 17460 12792
rect 17328 12406 17448 12434
rect 17316 12368 17368 12374
rect 17314 12336 17316 12345
rect 17368 12336 17370 12345
rect 17314 12271 17370 12280
rect 17224 10464 17276 10470
rect 17038 10432 17094 10441
rect 17224 10406 17276 10412
rect 16486 10364 16794 10373
rect 17038 10367 17094 10376
rect 16486 10362 16492 10364
rect 16548 10362 16572 10364
rect 16628 10362 16652 10364
rect 16708 10362 16732 10364
rect 16788 10362 16794 10364
rect 16548 10310 16550 10362
rect 16730 10310 16732 10362
rect 16486 10308 16492 10310
rect 16548 10308 16572 10310
rect 16628 10308 16652 10310
rect 16708 10308 16732 10310
rect 16788 10308 16794 10310
rect 16486 10299 16794 10308
rect 17052 10266 17080 10367
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 17420 10062 17448 12406
rect 17604 12374 17632 12872
rect 17776 12776 17828 12782
rect 17972 12730 18000 13670
rect 17776 12718 17828 12724
rect 17682 12608 17738 12617
rect 17682 12543 17738 12552
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17604 11150 17632 12310
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17696 10674 17724 12543
rect 17788 11830 17816 12718
rect 17880 12702 18000 12730
rect 17880 12442 17908 12702
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17972 10810 18000 12582
rect 18156 12322 18184 15830
rect 18248 15026 18276 16390
rect 18705 16348 19013 16357
rect 18705 16346 18711 16348
rect 18767 16346 18791 16348
rect 18847 16346 18871 16348
rect 18927 16346 18951 16348
rect 19007 16346 19013 16348
rect 18767 16294 18769 16346
rect 18949 16294 18951 16346
rect 18705 16292 18711 16294
rect 18767 16292 18791 16294
rect 18847 16292 18871 16294
rect 18927 16292 18951 16294
rect 19007 16292 19013 16294
rect 18705 16283 19013 16292
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18340 15026 18368 15506
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18248 13734 18276 14962
rect 18326 14920 18382 14929
rect 18326 14855 18382 14864
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18340 12434 18368 14855
rect 18432 13802 18460 15302
rect 18705 15260 19013 15269
rect 18705 15258 18711 15260
rect 18767 15258 18791 15260
rect 18847 15258 18871 15260
rect 18927 15258 18951 15260
rect 19007 15258 19013 15260
rect 18767 15206 18769 15258
rect 18949 15206 18951 15258
rect 18705 15204 18711 15206
rect 18767 15204 18791 15206
rect 18847 15204 18871 15206
rect 18927 15204 18951 15206
rect 19007 15204 19013 15206
rect 18705 15195 19013 15204
rect 19062 15056 19118 15065
rect 19118 15014 19196 15042
rect 19062 14991 19118 15000
rect 19062 14376 19118 14385
rect 19062 14311 19118 14320
rect 18705 14172 19013 14181
rect 18705 14170 18711 14172
rect 18767 14170 18791 14172
rect 18847 14170 18871 14172
rect 18927 14170 18951 14172
rect 19007 14170 19013 14172
rect 18767 14118 18769 14170
rect 18949 14118 18951 14170
rect 18705 14116 18711 14118
rect 18767 14116 18791 14118
rect 18847 14116 18871 14118
rect 18927 14116 18951 14118
rect 19007 14116 19013 14118
rect 18705 14107 19013 14116
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18510 13696 18566 13705
rect 18510 13631 18566 13640
rect 18064 12294 18184 12322
rect 18248 12406 18368 12434
rect 18418 12472 18474 12481
rect 18418 12407 18474 12416
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17512 10266 17540 10610
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17682 10024 17738 10033
rect 9827 9820 10135 9829
rect 9827 9818 9833 9820
rect 9889 9818 9913 9820
rect 9969 9818 9993 9820
rect 10049 9818 10073 9820
rect 10129 9818 10135 9820
rect 9889 9766 9891 9818
rect 10071 9766 10073 9818
rect 9827 9764 9833 9766
rect 9889 9764 9913 9766
rect 9969 9764 9993 9766
rect 10049 9764 10073 9766
rect 10129 9764 10135 9766
rect 9827 9755 10135 9764
rect 14266 9820 14574 9829
rect 14266 9818 14272 9820
rect 14328 9818 14352 9820
rect 14408 9818 14432 9820
rect 14488 9818 14512 9820
rect 14568 9818 14574 9820
rect 14328 9766 14330 9818
rect 14510 9766 14512 9818
rect 14266 9764 14272 9766
rect 14328 9764 14352 9766
rect 14408 9764 14432 9766
rect 14488 9764 14512 9766
rect 14568 9764 14574 9766
rect 14266 9755 14574 9764
rect 16960 9518 16988 9998
rect 17682 9959 17738 9968
rect 17696 9586 17724 9959
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 3169 9276 3477 9285
rect 3169 9274 3175 9276
rect 3231 9274 3255 9276
rect 3311 9274 3335 9276
rect 3391 9274 3415 9276
rect 3471 9274 3477 9276
rect 3231 9222 3233 9274
rect 3413 9222 3415 9274
rect 3169 9220 3175 9222
rect 3231 9220 3255 9222
rect 3311 9220 3335 9222
rect 3391 9220 3415 9222
rect 3471 9220 3477 9222
rect 3169 9211 3477 9220
rect 7608 9276 7916 9285
rect 7608 9274 7614 9276
rect 7670 9274 7694 9276
rect 7750 9274 7774 9276
rect 7830 9274 7854 9276
rect 7910 9274 7916 9276
rect 7670 9222 7672 9274
rect 7852 9222 7854 9274
rect 7608 9220 7614 9222
rect 7670 9220 7694 9222
rect 7750 9220 7774 9222
rect 7830 9220 7854 9222
rect 7910 9220 7916 9222
rect 7608 9211 7916 9220
rect 12047 9276 12355 9285
rect 12047 9274 12053 9276
rect 12109 9274 12133 9276
rect 12189 9274 12213 9276
rect 12269 9274 12293 9276
rect 12349 9274 12355 9276
rect 12109 9222 12111 9274
rect 12291 9222 12293 9274
rect 12047 9220 12053 9222
rect 12109 9220 12133 9222
rect 12189 9220 12213 9222
rect 12269 9220 12293 9222
rect 12349 9220 12355 9222
rect 12047 9211 12355 9220
rect 16486 9276 16794 9285
rect 16486 9274 16492 9276
rect 16548 9274 16572 9276
rect 16628 9274 16652 9276
rect 16708 9274 16732 9276
rect 16788 9274 16794 9276
rect 16548 9222 16550 9274
rect 16730 9222 16732 9274
rect 16486 9220 16492 9222
rect 16548 9220 16572 9222
rect 16628 9220 16652 9222
rect 16708 9220 16732 9222
rect 16788 9220 16794 9222
rect 16486 9211 16794 9220
rect 1584 8968 1636 8974
rect 1582 8936 1584 8945
rect 17040 8968 17092 8974
rect 1636 8936 1638 8945
rect 1582 8871 1638 8880
rect 17038 8936 17040 8945
rect 17092 8936 17094 8945
rect 17038 8871 17094 8880
rect 5388 8732 5696 8741
rect 5388 8730 5394 8732
rect 5450 8730 5474 8732
rect 5530 8730 5554 8732
rect 5610 8730 5634 8732
rect 5690 8730 5696 8732
rect 5450 8678 5452 8730
rect 5632 8678 5634 8730
rect 5388 8676 5394 8678
rect 5450 8676 5474 8678
rect 5530 8676 5554 8678
rect 5610 8676 5634 8678
rect 5690 8676 5696 8678
rect 5388 8667 5696 8676
rect 9827 8732 10135 8741
rect 9827 8730 9833 8732
rect 9889 8730 9913 8732
rect 9969 8730 9993 8732
rect 10049 8730 10073 8732
rect 10129 8730 10135 8732
rect 9889 8678 9891 8730
rect 10071 8678 10073 8730
rect 9827 8676 9833 8678
rect 9889 8676 9913 8678
rect 9969 8676 9993 8678
rect 10049 8676 10073 8678
rect 10129 8676 10135 8678
rect 9827 8667 10135 8676
rect 14266 8732 14574 8741
rect 14266 8730 14272 8732
rect 14328 8730 14352 8732
rect 14408 8730 14432 8732
rect 14488 8730 14512 8732
rect 14568 8730 14574 8732
rect 14328 8678 14330 8730
rect 14510 8678 14512 8730
rect 14266 8676 14272 8678
rect 14328 8676 14352 8678
rect 14408 8676 14432 8678
rect 14488 8676 14512 8678
rect 14568 8676 14574 8678
rect 14266 8667 14574 8676
rect 17038 8528 17094 8537
rect 18064 8498 18092 12294
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18156 11898 18184 12174
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18248 9178 18276 12406
rect 18326 11792 18382 11801
rect 18326 11727 18328 11736
rect 18380 11727 18382 11736
rect 18328 11698 18380 11704
rect 18326 11656 18382 11665
rect 18326 11591 18382 11600
rect 18340 11354 18368 11591
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18326 11248 18382 11257
rect 18326 11183 18382 11192
rect 18340 10266 18368 11183
rect 18432 10674 18460 12407
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18326 9208 18382 9217
rect 18236 9172 18288 9178
rect 18524 9178 18552 13631
rect 18705 13084 19013 13093
rect 18705 13082 18711 13084
rect 18767 13082 18791 13084
rect 18847 13082 18871 13084
rect 18927 13082 18951 13084
rect 19007 13082 19013 13084
rect 18767 13030 18769 13082
rect 18949 13030 18951 13082
rect 18705 13028 18711 13030
rect 18767 13028 18791 13030
rect 18847 13028 18871 13030
rect 18927 13028 18951 13030
rect 19007 13028 19013 13030
rect 18705 13019 19013 13028
rect 18705 11996 19013 12005
rect 18705 11994 18711 11996
rect 18767 11994 18791 11996
rect 18847 11994 18871 11996
rect 18927 11994 18951 11996
rect 19007 11994 19013 11996
rect 18767 11942 18769 11994
rect 18949 11942 18951 11994
rect 18705 11940 18711 11942
rect 18767 11940 18791 11942
rect 18847 11940 18871 11942
rect 18927 11940 18951 11942
rect 19007 11940 19013 11942
rect 18705 11931 19013 11940
rect 18705 10908 19013 10917
rect 18705 10906 18711 10908
rect 18767 10906 18791 10908
rect 18847 10906 18871 10908
rect 18927 10906 18951 10908
rect 19007 10906 19013 10908
rect 18767 10854 18769 10906
rect 18949 10854 18951 10906
rect 18705 10852 18711 10854
rect 18767 10852 18791 10854
rect 18847 10852 18871 10854
rect 18927 10852 18951 10854
rect 19007 10852 19013 10854
rect 18705 10843 19013 10852
rect 18602 10704 18658 10713
rect 18602 10639 18658 10648
rect 18616 9586 18644 10639
rect 18705 9820 19013 9829
rect 18705 9818 18711 9820
rect 18767 9818 18791 9820
rect 18847 9818 18871 9820
rect 18927 9818 18951 9820
rect 19007 9818 19013 9820
rect 18767 9766 18769 9818
rect 18949 9766 18951 9818
rect 18705 9764 18711 9766
rect 18767 9764 18791 9766
rect 18847 9764 18871 9766
rect 18927 9764 18951 9766
rect 19007 9764 19013 9766
rect 18705 9755 19013 9764
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18326 9143 18382 9152
rect 18512 9172 18564 9178
rect 18236 9114 18288 9120
rect 18340 8498 18368 9143
rect 18512 9114 18564 9120
rect 17038 8463 17040 8472
rect 17092 8463 17094 8472
rect 18052 8492 18104 8498
rect 17040 8434 17092 8440
rect 18052 8434 18104 8440
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 8129 1624 8298
rect 3169 8188 3477 8197
rect 3169 8186 3175 8188
rect 3231 8186 3255 8188
rect 3311 8186 3335 8188
rect 3391 8186 3415 8188
rect 3471 8186 3477 8188
rect 3231 8134 3233 8186
rect 3413 8134 3415 8186
rect 3169 8132 3175 8134
rect 3231 8132 3255 8134
rect 3311 8132 3335 8134
rect 3391 8132 3415 8134
rect 3471 8132 3477 8134
rect 1582 8120 1638 8129
rect 3169 8123 3477 8132
rect 7608 8188 7916 8197
rect 7608 8186 7614 8188
rect 7670 8186 7694 8188
rect 7750 8186 7774 8188
rect 7830 8186 7854 8188
rect 7910 8186 7916 8188
rect 7670 8134 7672 8186
rect 7852 8134 7854 8186
rect 7608 8132 7614 8134
rect 7670 8132 7694 8134
rect 7750 8132 7774 8134
rect 7830 8132 7854 8134
rect 7910 8132 7916 8134
rect 7608 8123 7916 8132
rect 12047 8188 12355 8197
rect 12047 8186 12053 8188
rect 12109 8186 12133 8188
rect 12189 8186 12213 8188
rect 12269 8186 12293 8188
rect 12349 8186 12355 8188
rect 12109 8134 12111 8186
rect 12291 8134 12293 8186
rect 12047 8132 12053 8134
rect 12109 8132 12133 8134
rect 12189 8132 12213 8134
rect 12269 8132 12293 8134
rect 12349 8132 12355 8134
rect 12047 8123 12355 8132
rect 16486 8188 16794 8197
rect 16486 8186 16492 8188
rect 16548 8186 16572 8188
rect 16628 8186 16652 8188
rect 16708 8186 16732 8188
rect 16788 8186 16794 8188
rect 16548 8134 16550 8186
rect 16730 8134 16732 8186
rect 16486 8132 16492 8134
rect 16548 8132 16572 8134
rect 16628 8132 16652 8134
rect 16708 8132 16732 8134
rect 16788 8132 16794 8134
rect 16486 8123 16794 8132
rect 18616 8090 18644 9522
rect 19076 9518 19104 14311
rect 19168 9654 19196 15014
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19260 9110 19288 19230
rect 19522 19200 19578 20000
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 18705 8732 19013 8741
rect 18705 8730 18711 8732
rect 18767 8730 18791 8732
rect 18847 8730 18871 8732
rect 18927 8730 18951 8732
rect 19007 8730 19013 8732
rect 18767 8678 18769 8730
rect 18949 8678 18951 8730
rect 18705 8676 18711 8678
rect 18767 8676 18791 8678
rect 18847 8676 18871 8678
rect 18927 8676 18951 8678
rect 19007 8676 19013 8678
rect 18705 8667 19013 8676
rect 1582 8055 1638 8064
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18326 7984 18382 7993
rect 18326 7919 18328 7928
rect 18380 7919 18382 7928
rect 18328 7890 18380 7896
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7721 1624 7822
rect 1582 7712 1638 7721
rect 1582 7647 1638 7656
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 18326 7440 18382 7449
rect 18326 7375 18328 7384
rect 18380 7375 18382 7384
rect 18328 7346 18380 7352
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6905 1624 7142
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1584 6792 1636 6798
rect 18328 6792 18380 6798
rect 1584 6734 1636 6740
rect 18326 6760 18328 6769
rect 18380 6760 18382 6769
rect 1596 6497 1624 6734
rect 18326 6695 18382 6704
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 1582 6488 1638 6497
rect 5388 6491 5696 6500
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 1582 6423 1638 6432
rect 18326 6352 18382 6361
rect 18326 6287 18328 6296
rect 18380 6287 18382 6296
rect 18328 6258 18380 6264
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 1584 5704 1636 5710
rect 1582 5672 1584 5681
rect 18328 5704 18380 5710
rect 1636 5672 1638 5681
rect 1582 5607 1638 5616
rect 18326 5672 18328 5681
rect 18380 5672 18382 5681
rect 18326 5607 18382 5616
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 1582 5264 1638 5273
rect 1582 5199 1584 5208
rect 1636 5199 1638 5208
rect 1584 5170 1636 5176
rect 18326 5128 18382 5137
rect 18326 5063 18328 5072
rect 18380 5063 18382 5072
rect 18328 5034 18380 5040
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 1596 4457 1624 4558
rect 1582 4448 1638 4457
rect 1582 4383 1638 4392
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 19168 4321 19196 4558
rect 19154 4312 19210 4321
rect 19154 4247 19210 4256
rect 1584 4072 1636 4078
rect 1582 4040 1584 4049
rect 1636 4040 1638 4049
rect 1582 3975 1638 3984
rect 18328 3936 18380 3942
rect 18326 3904 18328 3913
rect 18380 3904 18382 3913
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 16486 3836 16794 3845
rect 18326 3839 18382 3848
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 1596 3233 1624 3470
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 1582 3224 1638 3233
rect 5388 3227 5696 3236
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 1582 3159 1638 3168
rect 18340 3097 18368 3470
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 18326 3088 18382 3097
rect 18326 3023 18382 3032
rect 1584 2848 1636 2854
rect 1582 2816 1584 2825
rect 18328 2848 18380 2854
rect 1636 2816 1638 2825
rect 18328 2790 18380 2796
rect 1582 2751 1638 2760
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 18340 2689 18368 2790
rect 18326 2680 18382 2689
rect 18326 2615 18382 2624
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 1596 1601 1624 2382
rect 2240 2009 2268 2382
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 2226 2000 2282 2009
rect 2226 1935 2282 1944
rect 1582 1592 1638 1601
rect 1582 1527 1638 1536
rect 17696 1465 17724 2382
rect 18340 1873 18368 2382
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 18326 1864 18382 1873
rect 18326 1799 18382 1808
rect 17682 1456 17738 1465
rect 17682 1391 17738 1400
<< via2 >>
rect 2778 17856 2834 17912
rect 1398 16632 1454 16688
rect 1582 16224 1638 16280
rect 2870 17448 2926 17504
rect 3175 16890 3231 16892
rect 3255 16890 3311 16892
rect 3335 16890 3391 16892
rect 3415 16890 3471 16892
rect 3175 16838 3221 16890
rect 3221 16838 3231 16890
rect 3255 16838 3285 16890
rect 3285 16838 3297 16890
rect 3297 16838 3311 16890
rect 3335 16838 3349 16890
rect 3349 16838 3361 16890
rect 3361 16838 3391 16890
rect 3415 16838 3425 16890
rect 3425 16838 3471 16890
rect 3175 16836 3231 16838
rect 3255 16836 3311 16838
rect 3335 16836 3391 16838
rect 3415 16836 3471 16838
rect 5394 17434 5450 17436
rect 5474 17434 5530 17436
rect 5554 17434 5610 17436
rect 5634 17434 5690 17436
rect 5394 17382 5440 17434
rect 5440 17382 5450 17434
rect 5474 17382 5504 17434
rect 5504 17382 5516 17434
rect 5516 17382 5530 17434
rect 5554 17382 5568 17434
rect 5568 17382 5580 17434
rect 5580 17382 5610 17434
rect 5634 17382 5644 17434
rect 5644 17382 5690 17434
rect 5394 17380 5450 17382
rect 5474 17380 5530 17382
rect 5554 17380 5610 17382
rect 5634 17380 5690 17382
rect 5998 16516 6054 16552
rect 5998 16496 6000 16516
rect 6000 16496 6052 16516
rect 6052 16496 6054 16516
rect 5394 16346 5450 16348
rect 5474 16346 5530 16348
rect 5554 16346 5610 16348
rect 5634 16346 5690 16348
rect 5394 16294 5440 16346
rect 5440 16294 5450 16346
rect 5474 16294 5504 16346
rect 5504 16294 5516 16346
rect 5516 16294 5530 16346
rect 5554 16294 5568 16346
rect 5568 16294 5580 16346
rect 5580 16294 5610 16346
rect 5634 16294 5644 16346
rect 5644 16294 5690 16346
rect 5394 16292 5450 16294
rect 5474 16292 5530 16294
rect 5554 16292 5610 16294
rect 5634 16292 5690 16294
rect 5354 16108 5410 16144
rect 5354 16088 5356 16108
rect 5356 16088 5408 16108
rect 5408 16088 5410 16108
rect 3175 15802 3231 15804
rect 3255 15802 3311 15804
rect 3335 15802 3391 15804
rect 3415 15802 3471 15804
rect 3175 15750 3221 15802
rect 3221 15750 3231 15802
rect 3255 15750 3285 15802
rect 3285 15750 3297 15802
rect 3297 15750 3311 15802
rect 3335 15750 3349 15802
rect 3349 15750 3361 15802
rect 3361 15750 3391 15802
rect 3415 15750 3425 15802
rect 3425 15750 3471 15802
rect 3175 15748 3231 15750
rect 3255 15748 3311 15750
rect 3335 15748 3391 15750
rect 3415 15748 3471 15750
rect 1490 15408 1546 15464
rect 1582 15000 1638 15056
rect 3175 14714 3231 14716
rect 3255 14714 3311 14716
rect 3335 14714 3391 14716
rect 3415 14714 3471 14716
rect 3175 14662 3221 14714
rect 3221 14662 3231 14714
rect 3255 14662 3285 14714
rect 3285 14662 3297 14714
rect 3297 14662 3311 14714
rect 3335 14662 3349 14714
rect 3349 14662 3361 14714
rect 3361 14662 3391 14714
rect 3415 14662 3425 14714
rect 3425 14662 3471 14714
rect 3175 14660 3231 14662
rect 3255 14660 3311 14662
rect 3335 14660 3391 14662
rect 3415 14660 3471 14662
rect 1582 14184 1638 14240
rect 1582 13812 1584 13832
rect 1584 13812 1636 13832
rect 1636 13812 1638 13832
rect 1582 13776 1638 13812
rect 3175 13626 3231 13628
rect 3255 13626 3311 13628
rect 3335 13626 3391 13628
rect 3415 13626 3471 13628
rect 3175 13574 3221 13626
rect 3221 13574 3231 13626
rect 3255 13574 3285 13626
rect 3285 13574 3297 13626
rect 3297 13574 3311 13626
rect 3335 13574 3349 13626
rect 3349 13574 3361 13626
rect 3361 13574 3391 13626
rect 3415 13574 3425 13626
rect 3425 13574 3471 13626
rect 3175 13572 3231 13574
rect 3255 13572 3311 13574
rect 3335 13572 3391 13574
rect 3415 13572 3471 13574
rect 5394 15258 5450 15260
rect 5474 15258 5530 15260
rect 5554 15258 5610 15260
rect 5634 15258 5690 15260
rect 5394 15206 5440 15258
rect 5440 15206 5450 15258
rect 5474 15206 5504 15258
rect 5504 15206 5516 15258
rect 5516 15206 5530 15258
rect 5554 15206 5568 15258
rect 5568 15206 5580 15258
rect 5580 15206 5610 15258
rect 5634 15206 5644 15258
rect 5644 15206 5690 15258
rect 5394 15204 5450 15206
rect 5474 15204 5530 15206
rect 5554 15204 5610 15206
rect 5634 15204 5690 15206
rect 5394 14170 5450 14172
rect 5474 14170 5530 14172
rect 5554 14170 5610 14172
rect 5634 14170 5690 14172
rect 5394 14118 5440 14170
rect 5440 14118 5450 14170
rect 5474 14118 5504 14170
rect 5504 14118 5516 14170
rect 5516 14118 5530 14170
rect 5554 14118 5568 14170
rect 5568 14118 5580 14170
rect 5580 14118 5610 14170
rect 5634 14118 5644 14170
rect 5644 14118 5690 14170
rect 5394 14116 5450 14118
rect 5474 14116 5530 14118
rect 5554 14116 5610 14118
rect 5634 14116 5690 14118
rect 5262 13368 5318 13424
rect 5394 13082 5450 13084
rect 5474 13082 5530 13084
rect 5554 13082 5610 13084
rect 5634 13082 5690 13084
rect 5394 13030 5440 13082
rect 5440 13030 5450 13082
rect 5474 13030 5504 13082
rect 5504 13030 5516 13082
rect 5516 13030 5530 13082
rect 5554 13030 5568 13082
rect 5568 13030 5580 13082
rect 5580 13030 5610 13082
rect 5634 13030 5644 13082
rect 5644 13030 5690 13082
rect 5394 13028 5450 13030
rect 5474 13028 5530 13030
rect 5554 13028 5610 13030
rect 5634 13028 5690 13030
rect 1582 12960 1638 13016
rect 6826 15952 6882 16008
rect 1582 12588 1584 12608
rect 1584 12588 1636 12608
rect 1636 12588 1638 12608
rect 1582 12552 1638 12588
rect 3175 12538 3231 12540
rect 3255 12538 3311 12540
rect 3335 12538 3391 12540
rect 3415 12538 3471 12540
rect 3175 12486 3221 12538
rect 3221 12486 3231 12538
rect 3255 12486 3285 12538
rect 3285 12486 3297 12538
rect 3297 12486 3311 12538
rect 3335 12486 3349 12538
rect 3349 12486 3361 12538
rect 3361 12486 3391 12538
rect 3415 12486 3425 12538
rect 3425 12486 3471 12538
rect 3175 12484 3231 12486
rect 3255 12484 3311 12486
rect 3335 12484 3391 12486
rect 3415 12484 3471 12486
rect 5394 11994 5450 11996
rect 5474 11994 5530 11996
rect 5554 11994 5610 11996
rect 5634 11994 5690 11996
rect 5394 11942 5440 11994
rect 5440 11942 5450 11994
rect 5474 11942 5504 11994
rect 5504 11942 5516 11994
rect 5516 11942 5530 11994
rect 5554 11942 5568 11994
rect 5568 11942 5580 11994
rect 5580 11942 5610 11994
rect 5634 11942 5644 11994
rect 5644 11942 5690 11994
rect 5394 11940 5450 11942
rect 5474 11940 5530 11942
rect 5554 11940 5610 11942
rect 5634 11940 5690 11942
rect 1582 11736 1638 11792
rect 3175 11450 3231 11452
rect 3255 11450 3311 11452
rect 3335 11450 3391 11452
rect 3415 11450 3471 11452
rect 3175 11398 3221 11450
rect 3221 11398 3231 11450
rect 3255 11398 3285 11450
rect 3285 11398 3297 11450
rect 3297 11398 3311 11450
rect 3335 11398 3349 11450
rect 3349 11398 3361 11450
rect 3361 11398 3391 11450
rect 3415 11398 3425 11450
rect 3425 11398 3471 11450
rect 3175 11396 3231 11398
rect 3255 11396 3311 11398
rect 3335 11396 3391 11398
rect 3415 11396 3471 11398
rect 1582 11328 1638 11384
rect 5394 10906 5450 10908
rect 5474 10906 5530 10908
rect 5554 10906 5610 10908
rect 5634 10906 5690 10908
rect 5394 10854 5440 10906
rect 5440 10854 5450 10906
rect 5474 10854 5504 10906
rect 5504 10854 5516 10906
rect 5516 10854 5530 10906
rect 5554 10854 5568 10906
rect 5568 10854 5580 10906
rect 5580 10854 5610 10906
rect 5634 10854 5644 10906
rect 5644 10854 5690 10906
rect 5394 10852 5450 10854
rect 5474 10852 5530 10854
rect 5554 10852 5610 10854
rect 5634 10852 5690 10854
rect 1582 10548 1584 10568
rect 1584 10548 1636 10568
rect 1636 10548 1638 10568
rect 1582 10512 1638 10548
rect 3175 10362 3231 10364
rect 3255 10362 3311 10364
rect 3335 10362 3391 10364
rect 3415 10362 3471 10364
rect 3175 10310 3221 10362
rect 3221 10310 3231 10362
rect 3255 10310 3285 10362
rect 3285 10310 3297 10362
rect 3297 10310 3311 10362
rect 3335 10310 3349 10362
rect 3349 10310 3361 10362
rect 3361 10310 3391 10362
rect 3415 10310 3425 10362
rect 3425 10310 3471 10362
rect 3175 10308 3231 10310
rect 3255 10308 3311 10310
rect 3335 10308 3391 10310
rect 3415 10308 3471 10310
rect 1582 10140 1584 10160
rect 1584 10140 1636 10160
rect 1636 10140 1638 10160
rect 1582 10104 1638 10140
rect 5394 9818 5450 9820
rect 5474 9818 5530 9820
rect 5554 9818 5610 9820
rect 5634 9818 5690 9820
rect 5394 9766 5440 9818
rect 5440 9766 5450 9818
rect 5474 9766 5504 9818
rect 5504 9766 5516 9818
rect 5516 9766 5530 9818
rect 5554 9766 5568 9818
rect 5568 9766 5580 9818
rect 5580 9766 5610 9818
rect 5634 9766 5644 9818
rect 5644 9766 5690 9818
rect 5394 9764 5450 9766
rect 5474 9764 5530 9766
rect 5554 9764 5610 9766
rect 5634 9764 5690 9766
rect 7562 17176 7618 17232
rect 7378 17040 7434 17096
rect 8298 17212 8300 17232
rect 8300 17212 8352 17232
rect 8352 17212 8354 17232
rect 7614 16890 7670 16892
rect 7694 16890 7750 16892
rect 7774 16890 7830 16892
rect 7854 16890 7910 16892
rect 7614 16838 7660 16890
rect 7660 16838 7670 16890
rect 7694 16838 7724 16890
rect 7724 16838 7736 16890
rect 7736 16838 7750 16890
rect 7774 16838 7788 16890
rect 7788 16838 7800 16890
rect 7800 16838 7830 16890
rect 7854 16838 7864 16890
rect 7864 16838 7910 16890
rect 7614 16836 7670 16838
rect 7694 16836 7750 16838
rect 7774 16836 7830 16838
rect 7854 16836 7910 16838
rect 7746 15952 7802 16008
rect 7614 15802 7670 15804
rect 7694 15802 7750 15804
rect 7774 15802 7830 15804
rect 7854 15802 7910 15804
rect 7614 15750 7660 15802
rect 7660 15750 7670 15802
rect 7694 15750 7724 15802
rect 7724 15750 7736 15802
rect 7736 15750 7750 15802
rect 7774 15750 7788 15802
rect 7788 15750 7800 15802
rect 7800 15750 7830 15802
rect 7854 15750 7864 15802
rect 7864 15750 7910 15802
rect 7614 15748 7670 15750
rect 7694 15748 7750 15750
rect 7774 15748 7830 15750
rect 7854 15748 7910 15750
rect 8298 17176 8354 17212
rect 8574 17040 8630 17096
rect 7930 14864 7986 14920
rect 7614 14714 7670 14716
rect 7694 14714 7750 14716
rect 7774 14714 7830 14716
rect 7854 14714 7910 14716
rect 7614 14662 7660 14714
rect 7660 14662 7670 14714
rect 7694 14662 7724 14714
rect 7724 14662 7736 14714
rect 7736 14662 7750 14714
rect 7774 14662 7788 14714
rect 7788 14662 7800 14714
rect 7800 14662 7830 14714
rect 7854 14662 7864 14714
rect 7864 14662 7910 14714
rect 7614 14660 7670 14662
rect 7694 14660 7750 14662
rect 7774 14660 7830 14662
rect 7854 14660 7910 14662
rect 7614 13626 7670 13628
rect 7694 13626 7750 13628
rect 7774 13626 7830 13628
rect 7854 13626 7910 13628
rect 7614 13574 7660 13626
rect 7660 13574 7670 13626
rect 7694 13574 7724 13626
rect 7724 13574 7736 13626
rect 7736 13574 7750 13626
rect 7774 13574 7788 13626
rect 7788 13574 7800 13626
rect 7800 13574 7830 13626
rect 7854 13574 7864 13626
rect 7864 13574 7910 13626
rect 7614 13572 7670 13574
rect 7694 13572 7750 13574
rect 7774 13572 7830 13574
rect 7854 13572 7910 13574
rect 8298 16224 8354 16280
rect 8022 13232 8078 13288
rect 8666 15988 8668 16008
rect 8668 15988 8720 16008
rect 8720 15988 8722 16008
rect 8666 15952 8722 15988
rect 8942 15988 8944 16008
rect 8944 15988 8996 16008
rect 8996 15988 8998 16008
rect 8942 15952 8998 15988
rect 8758 15000 8814 15056
rect 7614 12538 7670 12540
rect 7694 12538 7750 12540
rect 7774 12538 7830 12540
rect 7854 12538 7910 12540
rect 7614 12486 7660 12538
rect 7660 12486 7670 12538
rect 7694 12486 7724 12538
rect 7724 12486 7736 12538
rect 7736 12486 7750 12538
rect 7774 12486 7788 12538
rect 7788 12486 7800 12538
rect 7800 12486 7830 12538
rect 7854 12486 7864 12538
rect 7864 12486 7910 12538
rect 7614 12484 7670 12486
rect 7694 12484 7750 12486
rect 7774 12484 7830 12486
rect 7854 12484 7910 12486
rect 9310 16088 9366 16144
rect 9833 17434 9889 17436
rect 9913 17434 9969 17436
rect 9993 17434 10049 17436
rect 10073 17434 10129 17436
rect 9833 17382 9879 17434
rect 9879 17382 9889 17434
rect 9913 17382 9943 17434
rect 9943 17382 9955 17434
rect 9955 17382 9969 17434
rect 9993 17382 10007 17434
rect 10007 17382 10019 17434
rect 10019 17382 10049 17434
rect 10073 17382 10083 17434
rect 10083 17382 10129 17434
rect 9833 17380 9889 17382
rect 9913 17380 9969 17382
rect 9993 17380 10049 17382
rect 10073 17380 10129 17382
rect 9494 16224 9550 16280
rect 10230 16788 10286 16824
rect 10230 16768 10232 16788
rect 10232 16768 10284 16788
rect 10284 16768 10286 16788
rect 9833 16346 9889 16348
rect 9913 16346 9969 16348
rect 9993 16346 10049 16348
rect 10073 16346 10129 16348
rect 9833 16294 9879 16346
rect 9879 16294 9889 16346
rect 9913 16294 9943 16346
rect 9943 16294 9955 16346
rect 9955 16294 9969 16346
rect 9993 16294 10007 16346
rect 10007 16294 10019 16346
rect 10019 16294 10049 16346
rect 10073 16294 10083 16346
rect 10083 16294 10129 16346
rect 9833 16292 9889 16294
rect 9913 16292 9969 16294
rect 9993 16292 10049 16294
rect 10073 16292 10129 16294
rect 9770 15580 9772 15600
rect 9772 15580 9824 15600
rect 9824 15580 9826 15600
rect 9770 15544 9826 15580
rect 9954 15408 10010 15464
rect 9494 14320 9550 14376
rect 9402 13932 9458 13968
rect 9402 13912 9404 13932
rect 9404 13912 9456 13932
rect 9456 13912 9458 13932
rect 9833 15258 9889 15260
rect 9913 15258 9969 15260
rect 9993 15258 10049 15260
rect 10073 15258 10129 15260
rect 9833 15206 9879 15258
rect 9879 15206 9889 15258
rect 9913 15206 9943 15258
rect 9943 15206 9955 15258
rect 9955 15206 9969 15258
rect 9993 15206 10007 15258
rect 10007 15206 10019 15258
rect 10019 15206 10049 15258
rect 10073 15206 10083 15258
rect 10083 15206 10129 15258
rect 9833 15204 9889 15206
rect 9913 15204 9969 15206
rect 9993 15204 10049 15206
rect 10073 15204 10129 15206
rect 10506 16224 10562 16280
rect 10138 14592 10194 14648
rect 9833 14170 9889 14172
rect 9913 14170 9969 14172
rect 9993 14170 10049 14172
rect 10073 14170 10129 14172
rect 9833 14118 9879 14170
rect 9879 14118 9889 14170
rect 9913 14118 9943 14170
rect 9943 14118 9955 14170
rect 9955 14118 9969 14170
rect 9993 14118 10007 14170
rect 10007 14118 10019 14170
rect 10019 14118 10049 14170
rect 10073 14118 10083 14170
rect 10083 14118 10129 14170
rect 9833 14116 9889 14118
rect 9913 14116 9969 14118
rect 9993 14116 10049 14118
rect 10073 14116 10129 14118
rect 10046 13776 10102 13832
rect 9833 13082 9889 13084
rect 9913 13082 9969 13084
rect 9993 13082 10049 13084
rect 10073 13082 10129 13084
rect 9833 13030 9879 13082
rect 9879 13030 9889 13082
rect 9913 13030 9943 13082
rect 9943 13030 9955 13082
rect 9955 13030 9969 13082
rect 9993 13030 10007 13082
rect 10007 13030 10019 13082
rect 10019 13030 10049 13082
rect 10073 13030 10083 13082
rect 10083 13030 10129 13082
rect 9833 13028 9889 13030
rect 9913 13028 9969 13030
rect 9993 13028 10049 13030
rect 10073 13028 10129 13030
rect 9833 11994 9889 11996
rect 9913 11994 9969 11996
rect 9993 11994 10049 11996
rect 10073 11994 10129 11996
rect 9833 11942 9879 11994
rect 9879 11942 9889 11994
rect 9913 11942 9943 11994
rect 9943 11942 9955 11994
rect 9955 11942 9969 11994
rect 9993 11942 10007 11994
rect 10007 11942 10019 11994
rect 10019 11942 10049 11994
rect 10073 11942 10083 11994
rect 10083 11942 10129 11994
rect 9833 11940 9889 11942
rect 9913 11940 9969 11942
rect 9993 11940 10049 11942
rect 10073 11940 10129 11942
rect 9126 11736 9182 11792
rect 10322 14456 10378 14512
rect 10598 15136 10654 15192
rect 10506 13676 10508 13696
rect 10508 13676 10560 13696
rect 10560 13676 10562 13696
rect 10506 13640 10562 13676
rect 10414 13504 10470 13560
rect 10506 12960 10562 13016
rect 10506 12844 10562 12880
rect 10506 12824 10508 12844
rect 10508 12824 10560 12844
rect 10560 12824 10562 12844
rect 10966 16768 11022 16824
rect 11058 16652 11114 16688
rect 11058 16632 11060 16652
rect 11060 16632 11112 16652
rect 11112 16632 11114 16652
rect 10874 14592 10930 14648
rect 10782 13640 10838 13696
rect 7614 11450 7670 11452
rect 7694 11450 7750 11452
rect 7774 11450 7830 11452
rect 7854 11450 7910 11452
rect 7614 11398 7660 11450
rect 7660 11398 7670 11450
rect 7694 11398 7724 11450
rect 7724 11398 7736 11450
rect 7736 11398 7750 11450
rect 7774 11398 7788 11450
rect 7788 11398 7800 11450
rect 7800 11398 7830 11450
rect 7854 11398 7864 11450
rect 7864 11398 7910 11450
rect 7614 11396 7670 11398
rect 7694 11396 7750 11398
rect 7774 11396 7830 11398
rect 7854 11396 7910 11398
rect 10690 12688 10746 12744
rect 15658 18944 15714 19000
rect 12053 16890 12109 16892
rect 12133 16890 12189 16892
rect 12213 16890 12269 16892
rect 12293 16890 12349 16892
rect 12053 16838 12099 16890
rect 12099 16838 12109 16890
rect 12133 16838 12163 16890
rect 12163 16838 12175 16890
rect 12175 16838 12189 16890
rect 12213 16838 12227 16890
rect 12227 16838 12239 16890
rect 12239 16838 12269 16890
rect 12293 16838 12303 16890
rect 12303 16838 12349 16890
rect 12053 16836 12109 16838
rect 12133 16836 12189 16838
rect 12213 16836 12269 16838
rect 12293 16836 12349 16838
rect 11058 15272 11114 15328
rect 11058 14184 11114 14240
rect 11242 14048 11298 14104
rect 11242 13812 11244 13832
rect 11244 13812 11296 13832
rect 11296 13812 11298 13832
rect 11242 13776 11298 13812
rect 11058 12844 11114 12880
rect 11058 12824 11060 12844
rect 11060 12824 11112 12844
rect 11112 12824 11114 12844
rect 11426 16360 11482 16416
rect 12254 16360 12310 16416
rect 12346 16224 12402 16280
rect 12053 15802 12109 15804
rect 12133 15802 12189 15804
rect 12213 15802 12269 15804
rect 12293 15802 12349 15804
rect 12053 15750 12099 15802
rect 12099 15750 12109 15802
rect 12133 15750 12163 15802
rect 12163 15750 12175 15802
rect 12175 15750 12189 15802
rect 12213 15750 12227 15802
rect 12227 15750 12239 15802
rect 12239 15750 12269 15802
rect 12293 15750 12303 15802
rect 12303 15750 12349 15802
rect 12053 15748 12109 15750
rect 12133 15748 12189 15750
rect 12213 15748 12269 15750
rect 12293 15748 12349 15750
rect 12714 15408 12770 15464
rect 11610 13776 11666 13832
rect 11610 13504 11666 13560
rect 11702 12280 11758 12336
rect 12053 14714 12109 14716
rect 12133 14714 12189 14716
rect 12213 14714 12269 14716
rect 12293 14714 12349 14716
rect 12053 14662 12099 14714
rect 12099 14662 12109 14714
rect 12133 14662 12163 14714
rect 12163 14662 12175 14714
rect 12175 14662 12189 14714
rect 12213 14662 12227 14714
rect 12227 14662 12239 14714
rect 12239 14662 12269 14714
rect 12293 14662 12303 14714
rect 12303 14662 12349 14714
rect 12053 14660 12109 14662
rect 12133 14660 12189 14662
rect 12213 14660 12269 14662
rect 12293 14660 12349 14662
rect 12254 14456 12310 14512
rect 12346 13776 12402 13832
rect 12530 13776 12586 13832
rect 12053 13626 12109 13628
rect 12133 13626 12189 13628
rect 12213 13626 12269 13628
rect 12293 13626 12349 13628
rect 12053 13574 12099 13626
rect 12099 13574 12109 13626
rect 12133 13574 12163 13626
rect 12163 13574 12175 13626
rect 12175 13574 12189 13626
rect 12213 13574 12227 13626
rect 12227 13574 12239 13626
rect 12239 13574 12269 13626
rect 12293 13574 12303 13626
rect 12303 13574 12349 13626
rect 12053 13572 12109 13574
rect 12133 13572 12189 13574
rect 12213 13572 12269 13574
rect 12293 13572 12349 13574
rect 12622 13504 12678 13560
rect 12162 12824 12218 12880
rect 14272 17434 14328 17436
rect 14352 17434 14408 17436
rect 14432 17434 14488 17436
rect 14512 17434 14568 17436
rect 14272 17382 14318 17434
rect 14318 17382 14328 17434
rect 14352 17382 14382 17434
rect 14382 17382 14394 17434
rect 14394 17382 14408 17434
rect 14432 17382 14446 17434
rect 14446 17382 14458 17434
rect 14458 17382 14488 17434
rect 14512 17382 14522 17434
rect 14522 17382 14568 17434
rect 14272 17380 14328 17382
rect 14352 17380 14408 17382
rect 14432 17380 14488 17382
rect 14512 17380 14568 17382
rect 13634 16632 13690 16688
rect 13174 15680 13230 15736
rect 13082 14456 13138 14512
rect 13082 14220 13084 14240
rect 13084 14220 13136 14240
rect 13136 14220 13138 14240
rect 13082 14184 13138 14220
rect 12898 13776 12954 13832
rect 12898 13640 12954 13696
rect 12053 12538 12109 12540
rect 12133 12538 12189 12540
rect 12213 12538 12269 12540
rect 12293 12538 12349 12540
rect 12053 12486 12099 12538
rect 12099 12486 12109 12538
rect 12133 12486 12163 12538
rect 12163 12486 12175 12538
rect 12175 12486 12189 12538
rect 12213 12486 12227 12538
rect 12227 12486 12239 12538
rect 12239 12486 12269 12538
rect 12293 12486 12303 12538
rect 12303 12486 12349 12538
rect 12053 12484 12109 12486
rect 12133 12484 12189 12486
rect 12213 12484 12269 12486
rect 12293 12484 12349 12486
rect 12622 12416 12678 12472
rect 13358 15816 13414 15872
rect 13266 14728 13322 14784
rect 13266 14456 13322 14512
rect 13358 13388 13414 13424
rect 13358 13368 13360 13388
rect 13360 13368 13412 13388
rect 13412 13368 13414 13388
rect 13358 12416 13414 12472
rect 13358 12280 13414 12336
rect 13450 11600 13506 11656
rect 12990 11464 13046 11520
rect 12053 11450 12109 11452
rect 12133 11450 12189 11452
rect 12213 11450 12269 11452
rect 12293 11450 12349 11452
rect 12053 11398 12099 11450
rect 12099 11398 12109 11450
rect 12133 11398 12163 11450
rect 12163 11398 12175 11450
rect 12175 11398 12189 11450
rect 12213 11398 12227 11450
rect 12227 11398 12239 11450
rect 12239 11398 12269 11450
rect 12293 11398 12303 11450
rect 12303 11398 12349 11450
rect 12053 11396 12109 11398
rect 12133 11396 12189 11398
rect 12213 11396 12269 11398
rect 12293 11396 12349 11398
rect 9833 10906 9889 10908
rect 9913 10906 9969 10908
rect 9993 10906 10049 10908
rect 10073 10906 10129 10908
rect 9833 10854 9879 10906
rect 9879 10854 9889 10906
rect 9913 10854 9943 10906
rect 9943 10854 9955 10906
rect 9955 10854 9969 10906
rect 9993 10854 10007 10906
rect 10007 10854 10019 10906
rect 10019 10854 10049 10906
rect 10073 10854 10083 10906
rect 10083 10854 10129 10906
rect 9833 10852 9889 10854
rect 9913 10852 9969 10854
rect 9993 10852 10049 10854
rect 10073 10852 10129 10854
rect 7614 10362 7670 10364
rect 7694 10362 7750 10364
rect 7774 10362 7830 10364
rect 7854 10362 7910 10364
rect 7614 10310 7660 10362
rect 7660 10310 7670 10362
rect 7694 10310 7724 10362
rect 7724 10310 7736 10362
rect 7736 10310 7750 10362
rect 7774 10310 7788 10362
rect 7788 10310 7800 10362
rect 7800 10310 7830 10362
rect 7854 10310 7864 10362
rect 7864 10310 7910 10362
rect 7614 10308 7670 10310
rect 7694 10308 7750 10310
rect 7774 10308 7830 10310
rect 7854 10308 7910 10310
rect 12053 10362 12109 10364
rect 12133 10362 12189 10364
rect 12213 10362 12269 10364
rect 12293 10362 12349 10364
rect 12053 10310 12099 10362
rect 12099 10310 12109 10362
rect 12133 10310 12163 10362
rect 12163 10310 12175 10362
rect 12175 10310 12189 10362
rect 12213 10310 12227 10362
rect 12227 10310 12239 10362
rect 12239 10310 12269 10362
rect 12293 10310 12303 10362
rect 12303 10310 12349 10362
rect 12053 10308 12109 10310
rect 12133 10308 12189 10310
rect 12213 10308 12269 10310
rect 12293 10308 12349 10310
rect 13818 15680 13874 15736
rect 14002 15136 14058 15192
rect 14646 17176 14702 17232
rect 14272 16346 14328 16348
rect 14352 16346 14408 16348
rect 14432 16346 14488 16348
rect 14512 16346 14568 16348
rect 14272 16294 14318 16346
rect 14318 16294 14328 16346
rect 14352 16294 14382 16346
rect 14382 16294 14394 16346
rect 14394 16294 14408 16346
rect 14432 16294 14446 16346
rect 14446 16294 14458 16346
rect 14458 16294 14488 16346
rect 14512 16294 14522 16346
rect 14522 16294 14568 16346
rect 14272 16292 14328 16294
rect 14352 16292 14408 16294
rect 14432 16292 14488 16294
rect 14512 16292 14568 16294
rect 14272 15258 14328 15260
rect 14352 15258 14408 15260
rect 14432 15258 14488 15260
rect 14512 15258 14568 15260
rect 14272 15206 14318 15258
rect 14318 15206 14328 15258
rect 14352 15206 14382 15258
rect 14382 15206 14394 15258
rect 14394 15206 14408 15258
rect 14432 15206 14446 15258
rect 14446 15206 14458 15258
rect 14458 15206 14488 15258
rect 14512 15206 14522 15258
rect 14522 15206 14568 15258
rect 14272 15204 14328 15206
rect 14352 15204 14408 15206
rect 14432 15204 14488 15206
rect 14512 15204 14568 15206
rect 13726 12280 13782 12336
rect 13818 11872 13874 11928
rect 14094 14728 14150 14784
rect 14002 13504 14058 13560
rect 14370 14728 14426 14784
rect 14738 14728 14794 14784
rect 14272 14170 14328 14172
rect 14352 14170 14408 14172
rect 14432 14170 14488 14172
rect 14512 14170 14568 14172
rect 14272 14118 14318 14170
rect 14318 14118 14328 14170
rect 14352 14118 14382 14170
rect 14382 14118 14394 14170
rect 14394 14118 14408 14170
rect 14432 14118 14446 14170
rect 14446 14118 14458 14170
rect 14458 14118 14488 14170
rect 14512 14118 14522 14170
rect 14522 14118 14568 14170
rect 14272 14116 14328 14118
rect 14352 14116 14408 14118
rect 14432 14116 14488 14118
rect 14512 14116 14568 14118
rect 14272 13082 14328 13084
rect 14352 13082 14408 13084
rect 14432 13082 14488 13084
rect 14512 13082 14568 13084
rect 14272 13030 14318 13082
rect 14318 13030 14328 13082
rect 14352 13030 14382 13082
rect 14382 13030 14394 13082
rect 14394 13030 14408 13082
rect 14432 13030 14446 13082
rect 14446 13030 14458 13082
rect 14458 13030 14488 13082
rect 14512 13030 14522 13082
rect 14522 13030 14568 13082
rect 14272 13028 14328 13030
rect 14352 13028 14408 13030
rect 14432 13028 14488 13030
rect 14512 13028 14568 13030
rect 14646 12824 14702 12880
rect 14002 12144 14058 12200
rect 14272 11994 14328 11996
rect 14352 11994 14408 11996
rect 14432 11994 14488 11996
rect 14512 11994 14568 11996
rect 14272 11942 14318 11994
rect 14318 11942 14328 11994
rect 14352 11942 14382 11994
rect 14382 11942 14394 11994
rect 14394 11942 14408 11994
rect 14432 11942 14446 11994
rect 14446 11942 14458 11994
rect 14458 11942 14488 11994
rect 14512 11942 14522 11994
rect 14522 11942 14568 11994
rect 14272 11940 14328 11942
rect 14352 11940 14408 11942
rect 14432 11940 14488 11942
rect 14512 11940 14568 11942
rect 14462 11464 14518 11520
rect 14278 11348 14334 11384
rect 14278 11328 14280 11348
rect 14280 11328 14332 11348
rect 14332 11328 14334 11348
rect 14272 10906 14328 10908
rect 14352 10906 14408 10908
rect 14432 10906 14488 10908
rect 14512 10906 14568 10908
rect 14272 10854 14318 10906
rect 14318 10854 14328 10906
rect 14352 10854 14382 10906
rect 14382 10854 14394 10906
rect 14394 10854 14408 10906
rect 14432 10854 14446 10906
rect 14446 10854 14458 10906
rect 14458 10854 14488 10906
rect 14512 10854 14522 10906
rect 14522 10854 14568 10906
rect 14272 10852 14328 10854
rect 14352 10852 14408 10854
rect 14432 10852 14488 10854
rect 14512 10852 14568 10854
rect 15014 15564 15070 15600
rect 15014 15544 15016 15564
rect 15016 15544 15068 15564
rect 15068 15544 15070 15564
rect 15198 15544 15254 15600
rect 15014 15272 15070 15328
rect 14922 14728 14978 14784
rect 15290 15272 15346 15328
rect 15198 14456 15254 14512
rect 15106 14320 15162 14376
rect 14922 14048 14978 14104
rect 14830 13368 14886 13424
rect 15014 13096 15070 13152
rect 15198 13640 15254 13696
rect 15106 12824 15162 12880
rect 14830 12144 14886 12200
rect 14922 12008 14978 12064
rect 15474 14592 15530 14648
rect 15842 16244 15898 16280
rect 15842 16224 15844 16244
rect 15844 16224 15896 16244
rect 15896 16224 15898 16244
rect 15658 14864 15714 14920
rect 15566 12180 15568 12200
rect 15568 12180 15620 12200
rect 15620 12180 15622 12200
rect 15566 12144 15622 12180
rect 15842 15408 15898 15464
rect 15842 13776 15898 13832
rect 15750 12008 15806 12064
rect 15750 11092 15752 11112
rect 15752 11092 15804 11112
rect 15804 11092 15806 11112
rect 15750 11056 15806 11092
rect 16026 17720 16082 17776
rect 16026 15000 16082 15056
rect 16492 16890 16548 16892
rect 16572 16890 16628 16892
rect 16652 16890 16708 16892
rect 16732 16890 16788 16892
rect 16492 16838 16538 16890
rect 16538 16838 16548 16890
rect 16572 16838 16602 16890
rect 16602 16838 16614 16890
rect 16614 16838 16628 16890
rect 16652 16838 16666 16890
rect 16666 16838 16678 16890
rect 16678 16838 16708 16890
rect 16732 16838 16742 16890
rect 16742 16838 16788 16890
rect 16492 16836 16548 16838
rect 16572 16836 16628 16838
rect 16652 16836 16708 16838
rect 16732 16836 16788 16838
rect 16854 16496 16910 16552
rect 16762 15952 16818 16008
rect 16302 15816 16358 15872
rect 16492 15802 16548 15804
rect 16572 15802 16628 15804
rect 16652 15802 16708 15804
rect 16732 15802 16788 15804
rect 16492 15750 16538 15802
rect 16538 15750 16548 15802
rect 16572 15750 16602 15802
rect 16602 15750 16614 15802
rect 16614 15750 16628 15802
rect 16652 15750 16666 15802
rect 16666 15750 16678 15802
rect 16678 15750 16708 15802
rect 16732 15750 16742 15802
rect 16742 15750 16788 15802
rect 16492 15748 16548 15750
rect 16572 15748 16628 15750
rect 16652 15748 16708 15750
rect 16732 15748 16788 15750
rect 16492 14714 16548 14716
rect 16572 14714 16628 14716
rect 16652 14714 16708 14716
rect 16732 14714 16788 14716
rect 16492 14662 16538 14714
rect 16538 14662 16548 14714
rect 16572 14662 16602 14714
rect 16602 14662 16614 14714
rect 16614 14662 16628 14714
rect 16652 14662 16666 14714
rect 16666 14662 16678 14714
rect 16678 14662 16708 14714
rect 16732 14662 16742 14714
rect 16742 14662 16788 14714
rect 16492 14660 16548 14662
rect 16572 14660 16628 14662
rect 16652 14660 16708 14662
rect 16732 14660 16788 14662
rect 16854 14456 16910 14512
rect 16492 13626 16548 13628
rect 16572 13626 16628 13628
rect 16652 13626 16708 13628
rect 16732 13626 16788 13628
rect 16492 13574 16538 13626
rect 16538 13574 16548 13626
rect 16572 13574 16602 13626
rect 16602 13574 16614 13626
rect 16614 13574 16628 13626
rect 16652 13574 16666 13626
rect 16666 13574 16678 13626
rect 16678 13574 16708 13626
rect 16732 13574 16742 13626
rect 16742 13574 16788 13626
rect 16492 13572 16548 13574
rect 16572 13572 16628 13574
rect 16652 13572 16708 13574
rect 16732 13572 16788 13574
rect 16670 13368 16726 13424
rect 16486 13232 16542 13288
rect 16762 13096 16818 13152
rect 16486 12824 16542 12880
rect 16118 12416 16174 12472
rect 16118 11736 16174 11792
rect 16578 12724 16580 12744
rect 16580 12724 16632 12744
rect 16632 12724 16634 12744
rect 16578 12688 16634 12724
rect 16492 12538 16548 12540
rect 16572 12538 16628 12540
rect 16652 12538 16708 12540
rect 16732 12538 16788 12540
rect 16492 12486 16538 12538
rect 16538 12486 16548 12538
rect 16572 12486 16602 12538
rect 16602 12486 16614 12538
rect 16614 12486 16628 12538
rect 16652 12486 16666 12538
rect 16666 12486 16678 12538
rect 16678 12486 16708 12538
rect 16732 12486 16742 12538
rect 16742 12486 16788 12538
rect 16492 12484 16548 12486
rect 16572 12484 16628 12486
rect 16652 12484 16708 12486
rect 16732 12484 16788 12486
rect 16762 11600 16818 11656
rect 16302 11464 16358 11520
rect 16492 11450 16548 11452
rect 16572 11450 16628 11452
rect 16652 11450 16708 11452
rect 16732 11450 16788 11452
rect 16492 11398 16538 11450
rect 16538 11398 16548 11450
rect 16572 11398 16602 11450
rect 16602 11398 16614 11450
rect 16614 11398 16628 11450
rect 16652 11398 16666 11450
rect 16666 11398 16678 11450
rect 16678 11398 16708 11450
rect 16732 11398 16742 11450
rect 16742 11398 16788 11450
rect 16492 11396 16548 11398
rect 16572 11396 16628 11398
rect 16652 11396 16708 11398
rect 16732 11396 16788 11398
rect 17314 15272 17370 15328
rect 18711 17434 18767 17436
rect 18791 17434 18847 17436
rect 18871 17434 18927 17436
rect 18951 17434 19007 17436
rect 18711 17382 18757 17434
rect 18757 17382 18767 17434
rect 18791 17382 18821 17434
rect 18821 17382 18833 17434
rect 18833 17382 18847 17434
rect 18871 17382 18885 17434
rect 18885 17382 18897 17434
rect 18897 17382 18927 17434
rect 18951 17382 18961 17434
rect 18961 17382 19007 17434
rect 18711 17380 18767 17382
rect 18791 17380 18847 17382
rect 18871 17380 18927 17382
rect 18951 17380 19007 17382
rect 19154 17312 19210 17368
rect 19062 17176 19118 17232
rect 17038 13232 17094 13288
rect 17222 13368 17278 13424
rect 17314 13232 17370 13288
rect 17222 12960 17278 13016
rect 17774 14048 17830 14104
rect 17682 12960 17738 13016
rect 18050 13912 18106 13968
rect 18050 13776 18106 13832
rect 17314 12316 17316 12336
rect 17316 12316 17368 12336
rect 17368 12316 17370 12336
rect 17314 12280 17370 12316
rect 17038 10376 17094 10432
rect 16492 10362 16548 10364
rect 16572 10362 16628 10364
rect 16652 10362 16708 10364
rect 16732 10362 16788 10364
rect 16492 10310 16538 10362
rect 16538 10310 16548 10362
rect 16572 10310 16602 10362
rect 16602 10310 16614 10362
rect 16614 10310 16628 10362
rect 16652 10310 16666 10362
rect 16666 10310 16678 10362
rect 16678 10310 16708 10362
rect 16732 10310 16742 10362
rect 16742 10310 16788 10362
rect 16492 10308 16548 10310
rect 16572 10308 16628 10310
rect 16652 10308 16708 10310
rect 16732 10308 16788 10310
rect 17682 12552 17738 12608
rect 18711 16346 18767 16348
rect 18791 16346 18847 16348
rect 18871 16346 18927 16348
rect 18951 16346 19007 16348
rect 18711 16294 18757 16346
rect 18757 16294 18767 16346
rect 18791 16294 18821 16346
rect 18821 16294 18833 16346
rect 18833 16294 18847 16346
rect 18871 16294 18885 16346
rect 18885 16294 18897 16346
rect 18897 16294 18927 16346
rect 18951 16294 18961 16346
rect 18961 16294 19007 16346
rect 18711 16292 18767 16294
rect 18791 16292 18847 16294
rect 18871 16292 18927 16294
rect 18951 16292 19007 16294
rect 18326 14864 18382 14920
rect 18711 15258 18767 15260
rect 18791 15258 18847 15260
rect 18871 15258 18927 15260
rect 18951 15258 19007 15260
rect 18711 15206 18757 15258
rect 18757 15206 18767 15258
rect 18791 15206 18821 15258
rect 18821 15206 18833 15258
rect 18833 15206 18847 15258
rect 18871 15206 18885 15258
rect 18885 15206 18897 15258
rect 18897 15206 18927 15258
rect 18951 15206 18961 15258
rect 18961 15206 19007 15258
rect 18711 15204 18767 15206
rect 18791 15204 18847 15206
rect 18871 15204 18927 15206
rect 18951 15204 19007 15206
rect 19062 15000 19118 15056
rect 19062 14320 19118 14376
rect 18711 14170 18767 14172
rect 18791 14170 18847 14172
rect 18871 14170 18927 14172
rect 18951 14170 19007 14172
rect 18711 14118 18757 14170
rect 18757 14118 18767 14170
rect 18791 14118 18821 14170
rect 18821 14118 18833 14170
rect 18833 14118 18847 14170
rect 18871 14118 18885 14170
rect 18885 14118 18897 14170
rect 18897 14118 18927 14170
rect 18951 14118 18961 14170
rect 18961 14118 19007 14170
rect 18711 14116 18767 14118
rect 18791 14116 18847 14118
rect 18871 14116 18927 14118
rect 18951 14116 19007 14118
rect 18510 13640 18566 13696
rect 18418 12416 18474 12472
rect 9833 9818 9889 9820
rect 9913 9818 9969 9820
rect 9993 9818 10049 9820
rect 10073 9818 10129 9820
rect 9833 9766 9879 9818
rect 9879 9766 9889 9818
rect 9913 9766 9943 9818
rect 9943 9766 9955 9818
rect 9955 9766 9969 9818
rect 9993 9766 10007 9818
rect 10007 9766 10019 9818
rect 10019 9766 10049 9818
rect 10073 9766 10083 9818
rect 10083 9766 10129 9818
rect 9833 9764 9889 9766
rect 9913 9764 9969 9766
rect 9993 9764 10049 9766
rect 10073 9764 10129 9766
rect 14272 9818 14328 9820
rect 14352 9818 14408 9820
rect 14432 9818 14488 9820
rect 14512 9818 14568 9820
rect 14272 9766 14318 9818
rect 14318 9766 14328 9818
rect 14352 9766 14382 9818
rect 14382 9766 14394 9818
rect 14394 9766 14408 9818
rect 14432 9766 14446 9818
rect 14446 9766 14458 9818
rect 14458 9766 14488 9818
rect 14512 9766 14522 9818
rect 14522 9766 14568 9818
rect 14272 9764 14328 9766
rect 14352 9764 14408 9766
rect 14432 9764 14488 9766
rect 14512 9764 14568 9766
rect 17682 9968 17738 10024
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 3175 9274 3231 9276
rect 3255 9274 3311 9276
rect 3335 9274 3391 9276
rect 3415 9274 3471 9276
rect 3175 9222 3221 9274
rect 3221 9222 3231 9274
rect 3255 9222 3285 9274
rect 3285 9222 3297 9274
rect 3297 9222 3311 9274
rect 3335 9222 3349 9274
rect 3349 9222 3361 9274
rect 3361 9222 3391 9274
rect 3415 9222 3425 9274
rect 3425 9222 3471 9274
rect 3175 9220 3231 9222
rect 3255 9220 3311 9222
rect 3335 9220 3391 9222
rect 3415 9220 3471 9222
rect 7614 9274 7670 9276
rect 7694 9274 7750 9276
rect 7774 9274 7830 9276
rect 7854 9274 7910 9276
rect 7614 9222 7660 9274
rect 7660 9222 7670 9274
rect 7694 9222 7724 9274
rect 7724 9222 7736 9274
rect 7736 9222 7750 9274
rect 7774 9222 7788 9274
rect 7788 9222 7800 9274
rect 7800 9222 7830 9274
rect 7854 9222 7864 9274
rect 7864 9222 7910 9274
rect 7614 9220 7670 9222
rect 7694 9220 7750 9222
rect 7774 9220 7830 9222
rect 7854 9220 7910 9222
rect 12053 9274 12109 9276
rect 12133 9274 12189 9276
rect 12213 9274 12269 9276
rect 12293 9274 12349 9276
rect 12053 9222 12099 9274
rect 12099 9222 12109 9274
rect 12133 9222 12163 9274
rect 12163 9222 12175 9274
rect 12175 9222 12189 9274
rect 12213 9222 12227 9274
rect 12227 9222 12239 9274
rect 12239 9222 12269 9274
rect 12293 9222 12303 9274
rect 12303 9222 12349 9274
rect 12053 9220 12109 9222
rect 12133 9220 12189 9222
rect 12213 9220 12269 9222
rect 12293 9220 12349 9222
rect 16492 9274 16548 9276
rect 16572 9274 16628 9276
rect 16652 9274 16708 9276
rect 16732 9274 16788 9276
rect 16492 9222 16538 9274
rect 16538 9222 16548 9274
rect 16572 9222 16602 9274
rect 16602 9222 16614 9274
rect 16614 9222 16628 9274
rect 16652 9222 16666 9274
rect 16666 9222 16678 9274
rect 16678 9222 16708 9274
rect 16732 9222 16742 9274
rect 16742 9222 16788 9274
rect 16492 9220 16548 9222
rect 16572 9220 16628 9222
rect 16652 9220 16708 9222
rect 16732 9220 16788 9222
rect 1582 8916 1584 8936
rect 1584 8916 1636 8936
rect 1636 8916 1638 8936
rect 1582 8880 1638 8916
rect 17038 8916 17040 8936
rect 17040 8916 17092 8936
rect 17092 8916 17094 8936
rect 17038 8880 17094 8916
rect 5394 8730 5450 8732
rect 5474 8730 5530 8732
rect 5554 8730 5610 8732
rect 5634 8730 5690 8732
rect 5394 8678 5440 8730
rect 5440 8678 5450 8730
rect 5474 8678 5504 8730
rect 5504 8678 5516 8730
rect 5516 8678 5530 8730
rect 5554 8678 5568 8730
rect 5568 8678 5580 8730
rect 5580 8678 5610 8730
rect 5634 8678 5644 8730
rect 5644 8678 5690 8730
rect 5394 8676 5450 8678
rect 5474 8676 5530 8678
rect 5554 8676 5610 8678
rect 5634 8676 5690 8678
rect 9833 8730 9889 8732
rect 9913 8730 9969 8732
rect 9993 8730 10049 8732
rect 10073 8730 10129 8732
rect 9833 8678 9879 8730
rect 9879 8678 9889 8730
rect 9913 8678 9943 8730
rect 9943 8678 9955 8730
rect 9955 8678 9969 8730
rect 9993 8678 10007 8730
rect 10007 8678 10019 8730
rect 10019 8678 10049 8730
rect 10073 8678 10083 8730
rect 10083 8678 10129 8730
rect 9833 8676 9889 8678
rect 9913 8676 9969 8678
rect 9993 8676 10049 8678
rect 10073 8676 10129 8678
rect 14272 8730 14328 8732
rect 14352 8730 14408 8732
rect 14432 8730 14488 8732
rect 14512 8730 14568 8732
rect 14272 8678 14318 8730
rect 14318 8678 14328 8730
rect 14352 8678 14382 8730
rect 14382 8678 14394 8730
rect 14394 8678 14408 8730
rect 14432 8678 14446 8730
rect 14446 8678 14458 8730
rect 14458 8678 14488 8730
rect 14512 8678 14522 8730
rect 14522 8678 14568 8730
rect 14272 8676 14328 8678
rect 14352 8676 14408 8678
rect 14432 8676 14488 8678
rect 14512 8676 14568 8678
rect 17038 8492 17094 8528
rect 18326 11756 18382 11792
rect 18326 11736 18328 11756
rect 18328 11736 18380 11756
rect 18380 11736 18382 11756
rect 18326 11600 18382 11656
rect 18326 11192 18382 11248
rect 18326 9152 18382 9208
rect 18711 13082 18767 13084
rect 18791 13082 18847 13084
rect 18871 13082 18927 13084
rect 18951 13082 19007 13084
rect 18711 13030 18757 13082
rect 18757 13030 18767 13082
rect 18791 13030 18821 13082
rect 18821 13030 18833 13082
rect 18833 13030 18847 13082
rect 18871 13030 18885 13082
rect 18885 13030 18897 13082
rect 18897 13030 18927 13082
rect 18951 13030 18961 13082
rect 18961 13030 19007 13082
rect 18711 13028 18767 13030
rect 18791 13028 18847 13030
rect 18871 13028 18927 13030
rect 18951 13028 19007 13030
rect 18711 11994 18767 11996
rect 18791 11994 18847 11996
rect 18871 11994 18927 11996
rect 18951 11994 19007 11996
rect 18711 11942 18757 11994
rect 18757 11942 18767 11994
rect 18791 11942 18821 11994
rect 18821 11942 18833 11994
rect 18833 11942 18847 11994
rect 18871 11942 18885 11994
rect 18885 11942 18897 11994
rect 18897 11942 18927 11994
rect 18951 11942 18961 11994
rect 18961 11942 19007 11994
rect 18711 11940 18767 11942
rect 18791 11940 18847 11942
rect 18871 11940 18927 11942
rect 18951 11940 19007 11942
rect 18711 10906 18767 10908
rect 18791 10906 18847 10908
rect 18871 10906 18927 10908
rect 18951 10906 19007 10908
rect 18711 10854 18757 10906
rect 18757 10854 18767 10906
rect 18791 10854 18821 10906
rect 18821 10854 18833 10906
rect 18833 10854 18847 10906
rect 18871 10854 18885 10906
rect 18885 10854 18897 10906
rect 18897 10854 18927 10906
rect 18951 10854 18961 10906
rect 18961 10854 19007 10906
rect 18711 10852 18767 10854
rect 18791 10852 18847 10854
rect 18871 10852 18927 10854
rect 18951 10852 19007 10854
rect 18602 10648 18658 10704
rect 18711 9818 18767 9820
rect 18791 9818 18847 9820
rect 18871 9818 18927 9820
rect 18951 9818 19007 9820
rect 18711 9766 18757 9818
rect 18757 9766 18767 9818
rect 18791 9766 18821 9818
rect 18821 9766 18833 9818
rect 18833 9766 18847 9818
rect 18871 9766 18885 9818
rect 18885 9766 18897 9818
rect 18897 9766 18927 9818
rect 18951 9766 18961 9818
rect 18961 9766 19007 9818
rect 18711 9764 18767 9766
rect 18791 9764 18847 9766
rect 18871 9764 18927 9766
rect 18951 9764 19007 9766
rect 17038 8472 17040 8492
rect 17040 8472 17092 8492
rect 17092 8472 17094 8492
rect 3175 8186 3231 8188
rect 3255 8186 3311 8188
rect 3335 8186 3391 8188
rect 3415 8186 3471 8188
rect 3175 8134 3221 8186
rect 3221 8134 3231 8186
rect 3255 8134 3285 8186
rect 3285 8134 3297 8186
rect 3297 8134 3311 8186
rect 3335 8134 3349 8186
rect 3349 8134 3361 8186
rect 3361 8134 3391 8186
rect 3415 8134 3425 8186
rect 3425 8134 3471 8186
rect 3175 8132 3231 8134
rect 3255 8132 3311 8134
rect 3335 8132 3391 8134
rect 3415 8132 3471 8134
rect 7614 8186 7670 8188
rect 7694 8186 7750 8188
rect 7774 8186 7830 8188
rect 7854 8186 7910 8188
rect 7614 8134 7660 8186
rect 7660 8134 7670 8186
rect 7694 8134 7724 8186
rect 7724 8134 7736 8186
rect 7736 8134 7750 8186
rect 7774 8134 7788 8186
rect 7788 8134 7800 8186
rect 7800 8134 7830 8186
rect 7854 8134 7864 8186
rect 7864 8134 7910 8186
rect 7614 8132 7670 8134
rect 7694 8132 7750 8134
rect 7774 8132 7830 8134
rect 7854 8132 7910 8134
rect 12053 8186 12109 8188
rect 12133 8186 12189 8188
rect 12213 8186 12269 8188
rect 12293 8186 12349 8188
rect 12053 8134 12099 8186
rect 12099 8134 12109 8186
rect 12133 8134 12163 8186
rect 12163 8134 12175 8186
rect 12175 8134 12189 8186
rect 12213 8134 12227 8186
rect 12227 8134 12239 8186
rect 12239 8134 12269 8186
rect 12293 8134 12303 8186
rect 12303 8134 12349 8186
rect 12053 8132 12109 8134
rect 12133 8132 12189 8134
rect 12213 8132 12269 8134
rect 12293 8132 12349 8134
rect 16492 8186 16548 8188
rect 16572 8186 16628 8188
rect 16652 8186 16708 8188
rect 16732 8186 16788 8188
rect 16492 8134 16538 8186
rect 16538 8134 16548 8186
rect 16572 8134 16602 8186
rect 16602 8134 16614 8186
rect 16614 8134 16628 8186
rect 16652 8134 16666 8186
rect 16666 8134 16678 8186
rect 16678 8134 16708 8186
rect 16732 8134 16742 8186
rect 16742 8134 16788 8186
rect 16492 8132 16548 8134
rect 16572 8132 16628 8134
rect 16652 8132 16708 8134
rect 16732 8132 16788 8134
rect 1582 8064 1638 8120
rect 18711 8730 18767 8732
rect 18791 8730 18847 8732
rect 18871 8730 18927 8732
rect 18951 8730 19007 8732
rect 18711 8678 18757 8730
rect 18757 8678 18767 8730
rect 18791 8678 18821 8730
rect 18821 8678 18833 8730
rect 18833 8678 18847 8730
rect 18871 8678 18885 8730
rect 18885 8678 18897 8730
rect 18897 8678 18927 8730
rect 18951 8678 18961 8730
rect 18961 8678 19007 8730
rect 18711 8676 18767 8678
rect 18791 8676 18847 8678
rect 18871 8676 18927 8678
rect 18951 8676 19007 8678
rect 18326 7948 18382 7984
rect 18326 7928 18328 7948
rect 18328 7928 18380 7948
rect 18380 7928 18382 7948
rect 1582 7656 1638 7712
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 18326 7404 18382 7440
rect 18326 7384 18328 7404
rect 18328 7384 18380 7404
rect 18380 7384 18382 7404
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 1582 6840 1638 6896
rect 18326 6740 18328 6760
rect 18328 6740 18380 6760
rect 18380 6740 18382 6760
rect 18326 6704 18382 6740
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 1582 6432 1638 6488
rect 18326 6316 18382 6352
rect 18326 6296 18328 6316
rect 18328 6296 18380 6316
rect 18380 6296 18382 6316
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 1582 5652 1584 5672
rect 1584 5652 1636 5672
rect 1636 5652 1638 5672
rect 1582 5616 1638 5652
rect 18326 5652 18328 5672
rect 18328 5652 18380 5672
rect 18380 5652 18382 5672
rect 18326 5616 18382 5652
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 1582 5228 1638 5264
rect 1582 5208 1584 5228
rect 1584 5208 1636 5228
rect 1636 5208 1638 5228
rect 18326 5092 18382 5128
rect 18326 5072 18328 5092
rect 18328 5072 18380 5092
rect 18380 5072 18382 5092
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 1582 4392 1638 4448
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 19154 4256 19210 4312
rect 1582 4020 1584 4040
rect 1584 4020 1636 4040
rect 1636 4020 1638 4040
rect 1582 3984 1638 4020
rect 18326 3884 18328 3904
rect 18328 3884 18380 3904
rect 18380 3884 18382 3904
rect 18326 3848 18382 3884
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 1582 3168 1638 3224
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 18326 3032 18382 3088
rect 1582 2796 1584 2816
rect 1584 2796 1636 2816
rect 1636 2796 1638 2816
rect 1582 2760 1638 2796
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 18326 2624 18382 2680
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 2226 1944 2282 2000
rect 1582 1536 1638 1592
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
rect 18326 1808 18382 1864
rect 17682 1400 17738 1456
<< metal3 >>
rect 15653 19002 15719 19005
rect 19200 19002 20000 19032
rect 15653 19000 20000 19002
rect 15653 18944 15658 19000
rect 15714 18944 20000 19000
rect 15653 18942 20000 18944
rect 15653 18939 15719 18942
rect 19200 18912 20000 18942
rect 16246 18532 16252 18596
rect 16316 18594 16322 18596
rect 19200 18594 20000 18624
rect 16316 18534 20000 18594
rect 16316 18532 16322 18534
rect 19200 18504 20000 18534
rect 0 18232 800 18352
rect 19200 18096 20000 18216
rect 0 17914 800 17944
rect 2773 17914 2839 17917
rect 0 17912 2839 17914
rect 0 17856 2778 17912
rect 2834 17856 2839 17912
rect 0 17854 2839 17856
rect 0 17824 800 17854
rect 2773 17851 2839 17854
rect 16021 17778 16087 17781
rect 19200 17778 20000 17808
rect 16021 17776 20000 17778
rect 16021 17720 16026 17776
rect 16082 17720 20000 17776
rect 16021 17718 20000 17720
rect 16021 17715 16087 17718
rect 19200 17688 20000 17718
rect 0 17506 800 17536
rect 2865 17506 2931 17509
rect 0 17504 2931 17506
rect 0 17448 2870 17504
rect 2926 17448 2931 17504
rect 0 17446 2931 17448
rect 0 17416 800 17446
rect 2865 17443 2931 17446
rect 5384 17440 5700 17441
rect 5384 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5700 17440
rect 5384 17375 5700 17376
rect 9823 17440 10139 17441
rect 9823 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10139 17440
rect 9823 17375 10139 17376
rect 14262 17440 14578 17441
rect 14262 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14578 17440
rect 14262 17375 14578 17376
rect 18701 17440 19017 17441
rect 18701 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19017 17440
rect 18701 17375 19017 17376
rect 19200 17373 20000 17400
rect 19149 17368 20000 17373
rect 19149 17312 19154 17368
rect 19210 17312 20000 17368
rect 19149 17307 20000 17312
rect 19200 17280 20000 17307
rect 7557 17234 7623 17237
rect 8293 17234 8359 17237
rect 7557 17232 8359 17234
rect 7557 17176 7562 17232
rect 7618 17176 8298 17232
rect 8354 17176 8359 17232
rect 7557 17174 8359 17176
rect 7557 17171 7623 17174
rect 8293 17171 8359 17174
rect 14641 17234 14707 17237
rect 19057 17234 19123 17237
rect 14641 17232 19123 17234
rect 14641 17176 14646 17232
rect 14702 17176 19062 17232
rect 19118 17176 19123 17232
rect 14641 17174 19123 17176
rect 14641 17171 14707 17174
rect 19057 17171 19123 17174
rect 0 17008 800 17128
rect 7373 17098 7439 17101
rect 8569 17098 8635 17101
rect 7373 17096 8635 17098
rect 7373 17040 7378 17096
rect 7434 17040 8574 17096
rect 8630 17040 8635 17096
rect 7373 17038 8635 17040
rect 7373 17035 7439 17038
rect 8569 17035 8635 17038
rect 3165 16896 3481 16897
rect 3165 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3481 16896
rect 3165 16831 3481 16832
rect 7604 16896 7920 16897
rect 7604 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7920 16896
rect 7604 16831 7920 16832
rect 12043 16896 12359 16897
rect 12043 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12359 16896
rect 12043 16831 12359 16832
rect 16482 16896 16798 16897
rect 16482 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16798 16896
rect 19200 16872 20000 16992
rect 16482 16831 16798 16832
rect 10225 16826 10291 16829
rect 10961 16826 11027 16829
rect 10225 16824 11027 16826
rect 10225 16768 10230 16824
rect 10286 16768 10966 16824
rect 11022 16768 11027 16824
rect 10225 16766 11027 16768
rect 10225 16763 10291 16766
rect 10961 16763 11027 16766
rect 0 16690 800 16720
rect 1393 16690 1459 16693
rect 0 16688 1459 16690
rect 0 16632 1398 16688
rect 1454 16632 1459 16688
rect 0 16630 1459 16632
rect 0 16600 800 16630
rect 1393 16627 1459 16630
rect 11053 16690 11119 16693
rect 13629 16690 13695 16693
rect 11053 16688 13695 16690
rect 11053 16632 11058 16688
rect 11114 16632 13634 16688
rect 13690 16632 13695 16688
rect 11053 16630 13695 16632
rect 11053 16627 11119 16630
rect 13629 16627 13695 16630
rect 5993 16554 6059 16557
rect 16849 16554 16915 16557
rect 19200 16554 20000 16584
rect 5993 16552 16915 16554
rect 5993 16496 5998 16552
rect 6054 16496 16854 16552
rect 16910 16496 16915 16552
rect 5993 16494 16915 16496
rect 5993 16491 6059 16494
rect 16849 16491 16915 16494
rect 16990 16494 20000 16554
rect 11421 16418 11487 16421
rect 12249 16418 12315 16421
rect 11421 16416 12315 16418
rect 11421 16360 11426 16416
rect 11482 16360 12254 16416
rect 12310 16360 12315 16416
rect 11421 16358 12315 16360
rect 11421 16355 11487 16358
rect 12249 16355 12315 16358
rect 5384 16352 5700 16353
rect 0 16282 800 16312
rect 5384 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5700 16352
rect 5384 16287 5700 16288
rect 9823 16352 10139 16353
rect 9823 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10139 16352
rect 9823 16287 10139 16288
rect 14262 16352 14578 16353
rect 14262 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14578 16352
rect 14262 16287 14578 16288
rect 1577 16282 1643 16285
rect 0 16280 1643 16282
rect 0 16224 1582 16280
rect 1638 16224 1643 16280
rect 0 16222 1643 16224
rect 0 16192 800 16222
rect 1577 16219 1643 16222
rect 8293 16282 8359 16285
rect 9489 16282 9555 16285
rect 8293 16280 9555 16282
rect 8293 16224 8298 16280
rect 8354 16224 9494 16280
rect 9550 16224 9555 16280
rect 8293 16222 9555 16224
rect 8293 16219 8359 16222
rect 9489 16219 9555 16222
rect 10501 16282 10567 16285
rect 12341 16282 12407 16285
rect 10501 16280 12407 16282
rect 10501 16224 10506 16280
rect 10562 16224 12346 16280
rect 12402 16224 12407 16280
rect 10501 16222 12407 16224
rect 10501 16219 10567 16222
rect 12341 16219 12407 16222
rect 15837 16284 15903 16285
rect 15837 16280 15884 16284
rect 15948 16282 15954 16284
rect 15837 16224 15842 16280
rect 15837 16220 15884 16224
rect 15948 16222 15994 16282
rect 15948 16220 15954 16222
rect 15837 16219 15903 16220
rect 5349 16146 5415 16149
rect 9305 16146 9371 16149
rect 5349 16144 9371 16146
rect 5349 16088 5354 16144
rect 5410 16088 9310 16144
rect 9366 16088 9371 16144
rect 5349 16086 9371 16088
rect 5349 16083 5415 16086
rect 9305 16083 9371 16086
rect 10542 16084 10548 16148
rect 10612 16146 10618 16148
rect 16990 16146 17050 16494
rect 19200 16464 20000 16494
rect 18701 16352 19017 16353
rect 18701 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19017 16352
rect 18701 16287 19017 16288
rect 19200 16146 20000 16176
rect 10612 16086 17050 16146
rect 17174 16086 20000 16146
rect 10612 16084 10618 16086
rect 6821 16010 6887 16013
rect 7741 16010 7807 16013
rect 8661 16010 8727 16013
rect 6821 16008 8727 16010
rect 6821 15952 6826 16008
rect 6882 15952 7746 16008
rect 7802 15952 8666 16008
rect 8722 15952 8727 16008
rect 6821 15950 8727 15952
rect 6821 15947 6887 15950
rect 7741 15947 7807 15950
rect 8661 15947 8727 15950
rect 8937 16010 9003 16013
rect 16757 16010 16823 16013
rect 8937 16008 16823 16010
rect 8937 15952 8942 16008
rect 8998 15952 16762 16008
rect 16818 15952 16823 16008
rect 8937 15950 16823 15952
rect 8937 15947 9003 15950
rect 16757 15947 16823 15950
rect 0 15784 800 15904
rect 13353 15874 13419 15877
rect 16297 15874 16363 15877
rect 13353 15872 16363 15874
rect 13353 15816 13358 15872
rect 13414 15816 16302 15872
rect 16358 15816 16363 15872
rect 13353 15814 16363 15816
rect 13353 15811 13419 15814
rect 16297 15811 16363 15814
rect 3165 15808 3481 15809
rect 3165 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3481 15808
rect 3165 15743 3481 15744
rect 7604 15808 7920 15809
rect 7604 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7920 15808
rect 7604 15743 7920 15744
rect 12043 15808 12359 15809
rect 12043 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12359 15808
rect 12043 15743 12359 15744
rect 16482 15808 16798 15809
rect 16482 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16798 15808
rect 16482 15743 16798 15744
rect 13169 15738 13235 15741
rect 13813 15738 13879 15741
rect 13169 15736 13879 15738
rect 13169 15680 13174 15736
rect 13230 15680 13818 15736
rect 13874 15680 13879 15736
rect 13169 15678 13879 15680
rect 13169 15675 13235 15678
rect 13813 15675 13879 15678
rect 9765 15602 9831 15605
rect 11094 15602 11100 15604
rect 9765 15600 11100 15602
rect 9765 15544 9770 15600
rect 9826 15544 11100 15600
rect 9765 15542 11100 15544
rect 9765 15539 9831 15542
rect 11094 15540 11100 15542
rect 11164 15602 11170 15604
rect 13854 15602 13860 15604
rect 11164 15542 13860 15602
rect 11164 15540 11170 15542
rect 13854 15540 13860 15542
rect 13924 15602 13930 15604
rect 15009 15602 15075 15605
rect 13924 15600 15075 15602
rect 13924 15544 15014 15600
rect 15070 15544 15075 15600
rect 13924 15542 15075 15544
rect 13924 15540 13930 15542
rect 15009 15539 15075 15542
rect 15193 15602 15259 15605
rect 17174 15602 17234 16086
rect 19200 16056 20000 16086
rect 19200 15648 20000 15768
rect 15193 15600 17234 15602
rect 15193 15544 15198 15600
rect 15254 15544 17234 15600
rect 15193 15542 17234 15544
rect 15193 15539 15259 15542
rect 0 15466 800 15496
rect 1485 15466 1551 15469
rect 0 15464 1551 15466
rect 0 15408 1490 15464
rect 1546 15408 1551 15464
rect 0 15406 1551 15408
rect 0 15376 800 15406
rect 1485 15403 1551 15406
rect 9949 15466 10015 15469
rect 12709 15466 12775 15469
rect 15837 15466 15903 15469
rect 9949 15464 10426 15466
rect 9949 15408 9954 15464
rect 10010 15408 10426 15464
rect 9949 15406 10426 15408
rect 9949 15403 10015 15406
rect 10366 15330 10426 15406
rect 12709 15464 15903 15466
rect 12709 15408 12714 15464
rect 12770 15408 15842 15464
rect 15898 15408 15903 15464
rect 12709 15406 15903 15408
rect 12709 15403 12775 15406
rect 15837 15403 15903 15406
rect 11053 15330 11119 15333
rect 10366 15328 11119 15330
rect 10366 15272 11058 15328
rect 11114 15272 11119 15328
rect 10366 15270 11119 15272
rect 11053 15267 11119 15270
rect 15009 15330 15075 15333
rect 15285 15330 15351 15333
rect 17309 15330 17375 15333
rect 19200 15330 20000 15360
rect 15009 15328 17375 15330
rect 15009 15272 15014 15328
rect 15070 15272 15290 15328
rect 15346 15272 17314 15328
rect 17370 15272 17375 15328
rect 15009 15270 17375 15272
rect 15009 15267 15075 15270
rect 15285 15267 15351 15270
rect 17309 15267 17375 15270
rect 5384 15264 5700 15265
rect 5384 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5700 15264
rect 5384 15199 5700 15200
rect 9823 15264 10139 15265
rect 9823 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10139 15264
rect 9823 15199 10139 15200
rect 14262 15264 14578 15265
rect 14262 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14578 15264
rect 14262 15199 14578 15200
rect 18701 15264 19017 15265
rect 18701 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19017 15264
rect 18701 15199 19017 15200
rect 19152 15240 20000 15330
rect 10593 15194 10659 15197
rect 13997 15194 14063 15197
rect 10593 15192 14063 15194
rect 10593 15136 10598 15192
rect 10654 15136 14002 15192
rect 14058 15136 14063 15192
rect 10593 15134 14063 15136
rect 10593 15131 10659 15134
rect 13997 15131 14063 15134
rect 19152 15092 19212 15240
rect 0 15058 800 15088
rect 19060 15061 19212 15092
rect 1577 15058 1643 15061
rect 0 15056 1643 15058
rect 0 15000 1582 15056
rect 1638 15000 1643 15056
rect 0 14998 1643 15000
rect 0 14968 800 14998
rect 1577 14995 1643 14998
rect 8753 15058 8819 15061
rect 16021 15058 16087 15061
rect 8753 15056 16087 15058
rect 8753 15000 8758 15056
rect 8814 15000 16026 15056
rect 16082 15000 16087 15056
rect 8753 14998 16087 15000
rect 8753 14995 8819 14998
rect 16021 14995 16087 14998
rect 19057 15056 19212 15061
rect 19057 15000 19062 15056
rect 19118 15032 19212 15056
rect 19118 15000 19123 15032
rect 19057 14995 19123 15000
rect 7925 14922 7991 14925
rect 15653 14922 15719 14925
rect 7925 14920 15719 14922
rect 7925 14864 7930 14920
rect 7986 14864 15658 14920
rect 15714 14864 15719 14920
rect 7925 14862 15719 14864
rect 7925 14859 7991 14862
rect 15653 14859 15719 14862
rect 18321 14922 18387 14925
rect 19200 14922 20000 14952
rect 18321 14920 20000 14922
rect 18321 14864 18326 14920
rect 18382 14864 20000 14920
rect 18321 14862 20000 14864
rect 18321 14859 18387 14862
rect 19200 14832 20000 14862
rect 13261 14786 13327 14789
rect 14089 14786 14155 14789
rect 13261 14784 14155 14786
rect 13261 14728 13266 14784
rect 13322 14728 14094 14784
rect 14150 14728 14155 14784
rect 13261 14726 14155 14728
rect 13261 14723 13327 14726
rect 14089 14723 14155 14726
rect 14365 14786 14431 14789
rect 14733 14786 14799 14789
rect 14917 14786 14983 14789
rect 14365 14784 14983 14786
rect 14365 14728 14370 14784
rect 14426 14728 14738 14784
rect 14794 14728 14922 14784
rect 14978 14728 14983 14784
rect 14365 14726 14983 14728
rect 14365 14723 14431 14726
rect 14733 14723 14799 14726
rect 14917 14723 14983 14726
rect 3165 14720 3481 14721
rect 0 14560 800 14680
rect 3165 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3481 14720
rect 3165 14655 3481 14656
rect 7604 14720 7920 14721
rect 7604 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7920 14720
rect 7604 14655 7920 14656
rect 12043 14720 12359 14721
rect 12043 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12359 14720
rect 12043 14655 12359 14656
rect 16482 14720 16798 14721
rect 16482 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16798 14720
rect 16482 14655 16798 14656
rect 10133 14650 10199 14653
rect 10869 14650 10935 14653
rect 15469 14650 15535 14653
rect 10133 14648 10935 14650
rect 10133 14592 10138 14648
rect 10194 14592 10874 14648
rect 10930 14592 10935 14648
rect 10133 14590 10935 14592
rect 10133 14587 10199 14590
rect 10869 14587 10935 14590
rect 12758 14648 15535 14650
rect 12758 14592 15474 14648
rect 15530 14592 15535 14648
rect 12758 14590 15535 14592
rect 10317 14514 10383 14517
rect 12249 14514 12315 14517
rect 12758 14514 12818 14590
rect 15469 14587 15535 14590
rect 10317 14512 12818 14514
rect 10317 14456 10322 14512
rect 10378 14456 12254 14512
rect 12310 14456 12818 14512
rect 10317 14454 12818 14456
rect 10317 14451 10383 14454
rect 12249 14451 12315 14454
rect 12934 14452 12940 14516
rect 13004 14514 13010 14516
rect 13077 14514 13143 14517
rect 13004 14512 13143 14514
rect 13004 14456 13082 14512
rect 13138 14456 13143 14512
rect 13004 14454 13143 14456
rect 13004 14452 13010 14454
rect 13077 14451 13143 14454
rect 13261 14514 13327 14517
rect 15193 14514 15259 14517
rect 13261 14512 15259 14514
rect 13261 14456 13266 14512
rect 13322 14456 15198 14512
rect 15254 14456 15259 14512
rect 13261 14454 15259 14456
rect 13261 14451 13327 14454
rect 15193 14451 15259 14454
rect 16062 14452 16068 14516
rect 16132 14514 16138 14516
rect 16849 14514 16915 14517
rect 16132 14512 16915 14514
rect 16132 14456 16854 14512
rect 16910 14456 16915 14512
rect 16132 14454 16915 14456
rect 16132 14452 16138 14454
rect 16849 14451 16915 14454
rect 19200 14424 20000 14544
rect 9489 14378 9555 14381
rect 15101 14378 15167 14381
rect 9489 14376 15167 14378
rect 9489 14320 9494 14376
rect 9550 14320 15106 14376
rect 15162 14320 15167 14376
rect 9489 14318 15167 14320
rect 9489 14315 9555 14318
rect 15101 14315 15167 14318
rect 19057 14376 19123 14381
rect 19057 14320 19062 14376
rect 19118 14344 19123 14376
rect 19118 14320 19212 14344
rect 19057 14315 19212 14320
rect 19060 14284 19212 14315
rect 0 14242 800 14272
rect 1577 14242 1643 14245
rect 0 14240 1643 14242
rect 0 14184 1582 14240
rect 1638 14184 1643 14240
rect 0 14182 1643 14184
rect 0 14152 800 14182
rect 1577 14179 1643 14182
rect 11053 14242 11119 14245
rect 13077 14242 13143 14245
rect 11053 14240 13143 14242
rect 11053 14184 11058 14240
rect 11114 14184 13082 14240
rect 13138 14184 13143 14240
rect 11053 14182 13143 14184
rect 11053 14179 11119 14182
rect 13077 14179 13143 14182
rect 5384 14176 5700 14177
rect 5384 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5700 14176
rect 5384 14111 5700 14112
rect 9823 14176 10139 14177
rect 9823 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10139 14176
rect 9823 14111 10139 14112
rect 14262 14176 14578 14177
rect 14262 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14578 14176
rect 14262 14111 14578 14112
rect 18701 14176 19017 14177
rect 18701 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19017 14176
rect 18701 14111 19017 14112
rect 19152 14136 19212 14284
rect 11094 14044 11100 14108
rect 11164 14106 11170 14108
rect 11237 14106 11303 14109
rect 11164 14104 11303 14106
rect 11164 14048 11242 14104
rect 11298 14048 11303 14104
rect 11164 14046 11303 14048
rect 11164 14044 11170 14046
rect 11237 14043 11303 14046
rect 14917 14106 14983 14109
rect 17769 14106 17835 14109
rect 14917 14104 17835 14106
rect 14917 14048 14922 14104
rect 14978 14048 17774 14104
rect 17830 14048 17835 14104
rect 14917 14046 17835 14048
rect 19152 14046 20000 14136
rect 14917 14043 14983 14046
rect 17769 14043 17835 14046
rect 19200 14016 20000 14046
rect 9397 13970 9463 13973
rect 18045 13970 18111 13973
rect 9397 13968 18111 13970
rect 9397 13912 9402 13968
rect 9458 13912 18050 13968
rect 18106 13912 18111 13968
rect 9397 13910 18111 13912
rect 9397 13907 9463 13910
rect 18045 13907 18111 13910
rect 0 13834 800 13864
rect 1577 13834 1643 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 800 13774
rect 1577 13771 1643 13774
rect 10041 13834 10107 13837
rect 11237 13834 11303 13837
rect 10041 13832 11303 13834
rect 10041 13776 10046 13832
rect 10102 13776 11242 13832
rect 11298 13776 11303 13832
rect 10041 13774 11303 13776
rect 10041 13771 10107 13774
rect 11237 13771 11303 13774
rect 11605 13834 11671 13837
rect 12341 13834 12407 13837
rect 11605 13832 12407 13834
rect 11605 13776 11610 13832
rect 11666 13776 12346 13832
rect 12402 13776 12407 13832
rect 11605 13774 12407 13776
rect 11605 13771 11671 13774
rect 12341 13771 12407 13774
rect 12525 13834 12591 13837
rect 12893 13834 12959 13837
rect 15694 13834 15700 13836
rect 12525 13832 15700 13834
rect 12525 13776 12530 13832
rect 12586 13776 12898 13832
rect 12954 13776 15700 13832
rect 12525 13774 15700 13776
rect 12525 13771 12591 13774
rect 12893 13771 12959 13774
rect 15694 13772 15700 13774
rect 15764 13834 15770 13836
rect 15837 13834 15903 13837
rect 18045 13834 18111 13837
rect 15764 13832 15903 13834
rect 15764 13776 15842 13832
rect 15898 13776 15903 13832
rect 15764 13774 15903 13776
rect 15764 13772 15770 13774
rect 15837 13771 15903 13774
rect 16300 13832 18111 13834
rect 16300 13776 18050 13832
rect 18106 13776 18111 13832
rect 16300 13774 18111 13776
rect 10501 13698 10567 13701
rect 10777 13698 10843 13701
rect 12893 13700 12959 13701
rect 12893 13698 12940 13700
rect 10501 13696 10843 13698
rect 10501 13640 10506 13696
rect 10562 13640 10782 13696
rect 10838 13640 10843 13696
rect 10501 13638 10843 13640
rect 12848 13696 12940 13698
rect 12848 13640 12898 13696
rect 12848 13638 12940 13640
rect 10501 13635 10567 13638
rect 10777 13635 10843 13638
rect 12893 13636 12940 13638
rect 13004 13636 13010 13700
rect 15193 13698 15259 13701
rect 16300 13698 16360 13774
rect 18045 13771 18111 13774
rect 15193 13696 16360 13698
rect 15193 13640 15198 13696
rect 15254 13640 16360 13696
rect 15193 13638 16360 13640
rect 18505 13698 18571 13701
rect 19200 13698 20000 13728
rect 18505 13696 20000 13698
rect 18505 13640 18510 13696
rect 18566 13640 20000 13696
rect 18505 13638 20000 13640
rect 12893 13635 12959 13636
rect 15193 13635 15259 13638
rect 18505 13635 18571 13638
rect 3165 13632 3481 13633
rect 3165 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3481 13632
rect 3165 13567 3481 13568
rect 7604 13632 7920 13633
rect 7604 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7920 13632
rect 7604 13567 7920 13568
rect 12043 13632 12359 13633
rect 12043 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12359 13632
rect 12043 13567 12359 13568
rect 16482 13632 16798 13633
rect 16482 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16798 13632
rect 19200 13608 20000 13638
rect 16482 13567 16798 13568
rect 10409 13562 10475 13565
rect 11605 13562 11671 13565
rect 10409 13560 11671 13562
rect 10409 13504 10414 13560
rect 10470 13504 11610 13560
rect 11666 13504 11671 13560
rect 10409 13502 11671 13504
rect 10409 13499 10475 13502
rect 11605 13499 11671 13502
rect 12617 13562 12683 13565
rect 13997 13562 14063 13565
rect 12617 13560 14063 13562
rect 12617 13504 12622 13560
rect 12678 13504 14002 13560
rect 14058 13504 14063 13560
rect 12617 13502 14063 13504
rect 12617 13499 12683 13502
rect 13997 13499 14063 13502
rect 0 13336 800 13456
rect 5257 13426 5323 13429
rect 13353 13426 13419 13429
rect 5257 13424 13419 13426
rect 5257 13368 5262 13424
rect 5318 13368 13358 13424
rect 13414 13368 13419 13424
rect 5257 13366 13419 13368
rect 5257 13363 5323 13366
rect 13353 13363 13419 13366
rect 14825 13426 14891 13429
rect 16665 13426 16731 13429
rect 17217 13426 17283 13429
rect 14825 13424 17283 13426
rect 14825 13368 14830 13424
rect 14886 13368 16670 13424
rect 16726 13368 17222 13424
rect 17278 13368 17283 13424
rect 14825 13366 17283 13368
rect 14825 13363 14891 13366
rect 16665 13363 16731 13366
rect 17217 13363 17283 13366
rect 8017 13290 8083 13293
rect 16481 13290 16547 13293
rect 17033 13292 17099 13293
rect 16982 13290 16988 13292
rect 8017 13288 16547 13290
rect 8017 13232 8022 13288
rect 8078 13232 16486 13288
rect 16542 13232 16547 13288
rect 8017 13230 16547 13232
rect 16942 13230 16988 13290
rect 17052 13288 17099 13292
rect 17094 13232 17099 13288
rect 8017 13227 8083 13230
rect 16481 13227 16547 13230
rect 16982 13228 16988 13230
rect 17052 13228 17099 13232
rect 17033 13227 17099 13228
rect 17309 13290 17375 13293
rect 19200 13290 20000 13320
rect 17309 13288 20000 13290
rect 17309 13232 17314 13288
rect 17370 13232 20000 13288
rect 17309 13230 20000 13232
rect 17309 13227 17375 13230
rect 19200 13200 20000 13230
rect 15009 13154 15075 13157
rect 16757 13154 16823 13157
rect 15009 13152 16823 13154
rect 15009 13096 15014 13152
rect 15070 13096 16762 13152
rect 16818 13096 16823 13152
rect 15009 13094 16823 13096
rect 15009 13091 15075 13094
rect 16757 13091 16823 13094
rect 5384 13088 5700 13089
rect 0 13018 800 13048
rect 5384 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5700 13088
rect 5384 13023 5700 13024
rect 9823 13088 10139 13089
rect 9823 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10139 13088
rect 9823 13023 10139 13024
rect 14262 13088 14578 13089
rect 14262 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14578 13088
rect 14262 13023 14578 13024
rect 18701 13088 19017 13089
rect 18701 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19017 13088
rect 18701 13023 19017 13024
rect 1577 13018 1643 13021
rect 0 13016 1643 13018
rect 0 12960 1582 13016
rect 1638 12960 1643 13016
rect 0 12958 1643 12960
rect 0 12928 800 12958
rect 1577 12955 1643 12958
rect 10501 13018 10567 13021
rect 17217 13018 17283 13021
rect 17677 13018 17743 13021
rect 10501 13016 14152 13018
rect 10501 12960 10506 13016
rect 10562 12960 14152 13016
rect 10501 12958 14152 12960
rect 10501 12955 10567 12958
rect 10501 12884 10567 12885
rect 10501 12882 10548 12884
rect 10456 12880 10548 12882
rect 10456 12824 10506 12880
rect 10456 12822 10548 12824
rect 10501 12820 10548 12822
rect 10612 12820 10618 12884
rect 11053 12882 11119 12885
rect 12157 12882 12223 12885
rect 11053 12880 12223 12882
rect 11053 12824 11058 12880
rect 11114 12824 12162 12880
rect 12218 12824 12223 12880
rect 11053 12822 12223 12824
rect 14092 12882 14152 12958
rect 17217 13016 17743 13018
rect 17217 12960 17222 13016
rect 17278 12960 17682 13016
rect 17738 12960 17743 13016
rect 17217 12958 17743 12960
rect 17217 12955 17283 12958
rect 17677 12955 17743 12958
rect 14641 12882 14707 12885
rect 15101 12882 15167 12885
rect 16481 12882 16547 12885
rect 19200 12882 20000 12912
rect 14092 12880 15167 12882
rect 14092 12824 14646 12880
rect 14702 12824 15106 12880
rect 15162 12824 15167 12880
rect 14092 12822 15167 12824
rect 10501 12819 10567 12820
rect 11053 12819 11119 12822
rect 12157 12819 12223 12822
rect 14641 12819 14707 12822
rect 15101 12819 15167 12822
rect 16116 12880 16547 12882
rect 16116 12824 16486 12880
rect 16542 12824 16547 12880
rect 16116 12822 16547 12824
rect 10685 12746 10751 12749
rect 16116 12746 16176 12822
rect 16481 12819 16547 12822
rect 17726 12822 20000 12882
rect 16573 12746 16639 12749
rect 10685 12744 16176 12746
rect 10685 12688 10690 12744
rect 10746 12688 16176 12744
rect 10685 12686 16176 12688
rect 16254 12744 16639 12746
rect 16254 12688 16578 12744
rect 16634 12688 16639 12744
rect 16254 12686 16639 12688
rect 10685 12683 10751 12686
rect 0 12610 800 12640
rect 1577 12610 1643 12613
rect 16254 12610 16314 12686
rect 16573 12683 16639 12686
rect 17726 12613 17786 12822
rect 19200 12792 20000 12822
rect 0 12608 1643 12610
rect 0 12552 1582 12608
rect 1638 12552 1643 12608
rect 0 12550 1643 12552
rect 0 12520 800 12550
rect 1577 12547 1643 12550
rect 12436 12550 16314 12610
rect 17677 12608 17786 12613
rect 17677 12552 17682 12608
rect 17738 12552 17786 12608
rect 17677 12550 17786 12552
rect 3165 12544 3481 12545
rect 3165 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3481 12544
rect 3165 12479 3481 12480
rect 7604 12544 7920 12545
rect 7604 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7920 12544
rect 7604 12479 7920 12480
rect 12043 12544 12359 12545
rect 12043 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12359 12544
rect 12043 12479 12359 12480
rect 11697 12338 11763 12341
rect 12436 12338 12496 12550
rect 17677 12547 17743 12550
rect 16482 12544 16798 12545
rect 16482 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16798 12544
rect 16482 12479 16798 12480
rect 12617 12474 12683 12477
rect 13353 12474 13419 12477
rect 16113 12476 16179 12477
rect 12617 12472 13419 12474
rect 12617 12416 12622 12472
rect 12678 12416 13358 12472
rect 13414 12416 13419 12472
rect 12617 12414 13419 12416
rect 12617 12411 12683 12414
rect 13353 12411 13419 12414
rect 16062 12412 16068 12476
rect 16132 12474 16179 12476
rect 18413 12474 18479 12477
rect 19200 12474 20000 12504
rect 16132 12472 16224 12474
rect 16174 12416 16224 12472
rect 16132 12414 16224 12416
rect 18413 12472 20000 12474
rect 18413 12416 18418 12472
rect 18474 12416 20000 12472
rect 18413 12414 20000 12416
rect 16132 12412 16179 12414
rect 16113 12411 16179 12412
rect 18413 12411 18479 12414
rect 19200 12384 20000 12414
rect 11697 12336 12496 12338
rect 11697 12280 11702 12336
rect 11758 12280 12496 12336
rect 11697 12278 12496 12280
rect 13353 12338 13419 12341
rect 13721 12338 13787 12341
rect 17309 12338 17375 12341
rect 13353 12336 17375 12338
rect 13353 12280 13358 12336
rect 13414 12280 13726 12336
rect 13782 12280 17314 12336
rect 17370 12280 17375 12336
rect 13353 12278 17375 12280
rect 11697 12275 11763 12278
rect 13353 12275 13419 12278
rect 13721 12275 13787 12278
rect 17309 12275 17375 12278
rect 0 12112 800 12232
rect 13997 12202 14063 12205
rect 14825 12202 14891 12205
rect 15561 12202 15627 12205
rect 13997 12200 14704 12202
rect 13997 12144 14002 12200
rect 14058 12144 14704 12200
rect 13997 12142 14704 12144
rect 13997 12139 14063 12142
rect 14644 12066 14704 12142
rect 14825 12200 15627 12202
rect 14825 12144 14830 12200
rect 14886 12144 15566 12200
rect 15622 12144 15627 12200
rect 14825 12142 15627 12144
rect 14825 12139 14891 12142
rect 15561 12139 15627 12142
rect 14917 12066 14983 12069
rect 14644 12064 14983 12066
rect 14644 12008 14922 12064
rect 14978 12008 14983 12064
rect 14644 12006 14983 12008
rect 14917 12003 14983 12006
rect 15745 12066 15811 12069
rect 15878 12066 15884 12068
rect 15745 12064 15884 12066
rect 15745 12008 15750 12064
rect 15806 12008 15884 12064
rect 15745 12006 15884 12008
rect 15745 12003 15811 12006
rect 15878 12004 15884 12006
rect 15948 12004 15954 12068
rect 19200 12066 20000 12096
rect 5384 12000 5700 12001
rect 5384 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5700 12000
rect 5384 11935 5700 11936
rect 9823 12000 10139 12001
rect 9823 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10139 12000
rect 9823 11935 10139 11936
rect 14262 12000 14578 12001
rect 14262 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14578 12000
rect 14262 11935 14578 11936
rect 18701 12000 19017 12001
rect 18701 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19017 12000
rect 18701 11935 19017 11936
rect 19152 11976 20000 12066
rect 13813 11932 13879 11933
rect 13813 11930 13860 11932
rect 13768 11928 13860 11930
rect 13768 11872 13818 11928
rect 13768 11870 13860 11872
rect 13813 11868 13860 11870
rect 13924 11868 13930 11932
rect 13813 11867 13879 11868
rect 19152 11828 19212 11976
rect 0 11794 800 11824
rect 1577 11794 1643 11797
rect 0 11792 1643 11794
rect 0 11736 1582 11792
rect 1638 11736 1643 11792
rect 0 11734 1643 11736
rect 0 11704 800 11734
rect 1577 11731 1643 11734
rect 9121 11794 9187 11797
rect 16113 11794 16179 11797
rect 9121 11792 16179 11794
rect 9121 11736 9126 11792
rect 9182 11736 16118 11792
rect 16174 11736 16179 11792
rect 9121 11734 16179 11736
rect 9121 11731 9187 11734
rect 16113 11731 16179 11734
rect 18321 11794 18387 11797
rect 19060 11794 19212 11828
rect 18321 11792 19212 11794
rect 18321 11736 18326 11792
rect 18382 11768 19212 11792
rect 18382 11736 19120 11768
rect 18321 11734 19120 11736
rect 18321 11731 18387 11734
rect 13445 11658 13511 11661
rect 16757 11658 16823 11661
rect 13445 11656 16823 11658
rect 13445 11600 13450 11656
rect 13506 11600 16762 11656
rect 16818 11600 16823 11656
rect 13445 11598 16823 11600
rect 13445 11595 13511 11598
rect 16757 11595 16823 11598
rect 18321 11658 18387 11661
rect 19200 11658 20000 11688
rect 18321 11656 20000 11658
rect 18321 11600 18326 11656
rect 18382 11600 20000 11656
rect 18321 11598 20000 11600
rect 18321 11595 18387 11598
rect 19200 11568 20000 11598
rect 12985 11522 13051 11525
rect 14457 11522 14523 11525
rect 16297 11522 16363 11525
rect 12985 11520 16363 11522
rect 12985 11464 12990 11520
rect 13046 11464 14462 11520
rect 14518 11464 16302 11520
rect 16358 11464 16363 11520
rect 12985 11462 16363 11464
rect 12985 11459 13051 11462
rect 14457 11459 14523 11462
rect 16297 11459 16363 11462
rect 3165 11456 3481 11457
rect 0 11386 800 11416
rect 3165 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3481 11456
rect 3165 11391 3481 11392
rect 7604 11456 7920 11457
rect 7604 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7920 11456
rect 7604 11391 7920 11392
rect 12043 11456 12359 11457
rect 12043 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12359 11456
rect 12043 11391 12359 11392
rect 16482 11456 16798 11457
rect 16482 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16798 11456
rect 16482 11391 16798 11392
rect 1577 11386 1643 11389
rect 0 11384 1643 11386
rect 0 11328 1582 11384
rect 1638 11328 1643 11384
rect 0 11326 1643 11328
rect 0 11296 800 11326
rect 1577 11323 1643 11326
rect 14273 11386 14339 11389
rect 15694 11386 15700 11388
rect 14273 11384 15700 11386
rect 14273 11328 14278 11384
rect 14334 11328 15700 11384
rect 14273 11326 15700 11328
rect 14273 11323 14339 11326
rect 15694 11324 15700 11326
rect 15764 11324 15770 11388
rect 18321 11250 18387 11253
rect 19200 11250 20000 11280
rect 18321 11248 20000 11250
rect 18321 11192 18326 11248
rect 18382 11192 20000 11248
rect 18321 11190 20000 11192
rect 18321 11187 18387 11190
rect 19200 11160 20000 11190
rect 15745 11114 15811 11117
rect 16982 11114 16988 11116
rect 15745 11112 16988 11114
rect 15745 11056 15750 11112
rect 15806 11056 16988 11112
rect 15745 11054 16988 11056
rect 15745 11051 15811 11054
rect 16982 11052 16988 11054
rect 17052 11052 17058 11116
rect 0 10888 800 11008
rect 5384 10912 5700 10913
rect 5384 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5700 10912
rect 5384 10847 5700 10848
rect 9823 10912 10139 10913
rect 9823 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10139 10912
rect 9823 10847 10139 10848
rect 14262 10912 14578 10913
rect 14262 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14578 10912
rect 14262 10847 14578 10848
rect 18701 10912 19017 10913
rect 18701 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19017 10912
rect 18701 10847 19017 10848
rect 19200 10842 20000 10872
rect 19152 10752 20000 10842
rect 18597 10706 18663 10709
rect 19152 10706 19212 10752
rect 18597 10704 19212 10706
rect 18597 10648 18602 10704
rect 18658 10648 19212 10704
rect 18597 10646 19212 10648
rect 18597 10643 18663 10646
rect 0 10570 800 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 800 10510
rect 1577 10507 1643 10510
rect 17033 10434 17099 10437
rect 19200 10434 20000 10464
rect 17033 10432 20000 10434
rect 17033 10376 17038 10432
rect 17094 10376 20000 10432
rect 17033 10374 20000 10376
rect 17033 10371 17099 10374
rect 3165 10368 3481 10369
rect 3165 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3481 10368
rect 3165 10303 3481 10304
rect 7604 10368 7920 10369
rect 7604 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7920 10368
rect 7604 10303 7920 10304
rect 12043 10368 12359 10369
rect 12043 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12359 10368
rect 12043 10303 12359 10304
rect 16482 10368 16798 10369
rect 16482 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16798 10368
rect 19200 10344 20000 10374
rect 16482 10303 16798 10304
rect 0 10162 800 10192
rect 1577 10162 1643 10165
rect 0 10160 1643 10162
rect 0 10104 1582 10160
rect 1638 10104 1643 10160
rect 0 10102 1643 10104
rect 0 10072 800 10102
rect 1577 10099 1643 10102
rect 17677 10026 17743 10029
rect 19200 10026 20000 10056
rect 17677 10024 20000 10026
rect 17677 9968 17682 10024
rect 17738 9968 20000 10024
rect 17677 9966 20000 9968
rect 17677 9963 17743 9966
rect 19200 9936 20000 9966
rect 5384 9824 5700 9825
rect 0 9664 800 9784
rect 5384 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5700 9824
rect 5384 9759 5700 9760
rect 9823 9824 10139 9825
rect 9823 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10139 9824
rect 9823 9759 10139 9760
rect 14262 9824 14578 9825
rect 14262 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14578 9824
rect 14262 9759 14578 9760
rect 18701 9824 19017 9825
rect 18701 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19017 9824
rect 18701 9759 19017 9760
rect 19200 9528 20000 9648
rect 0 9346 800 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 800 9286
rect 1577 9283 1643 9286
rect 3165 9280 3481 9281
rect 3165 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3481 9280
rect 3165 9215 3481 9216
rect 7604 9280 7920 9281
rect 7604 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7920 9280
rect 7604 9215 7920 9216
rect 12043 9280 12359 9281
rect 12043 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12359 9280
rect 12043 9215 12359 9216
rect 16482 9280 16798 9281
rect 16482 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16798 9280
rect 16482 9215 16798 9216
rect 18321 9210 18387 9213
rect 19200 9210 20000 9240
rect 18321 9208 20000 9210
rect 18321 9152 18326 9208
rect 18382 9152 20000 9208
rect 18321 9150 20000 9152
rect 18321 9147 18387 9150
rect 19200 9120 20000 9150
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 17033 8938 17099 8941
rect 17033 8936 19212 8938
rect 17033 8880 17038 8936
rect 17094 8880 19212 8936
rect 17033 8878 19212 8880
rect 17033 8875 17099 8878
rect 19152 8832 19212 8878
rect 19152 8742 20000 8832
rect 5384 8736 5700 8737
rect 5384 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5700 8736
rect 5384 8671 5700 8672
rect 9823 8736 10139 8737
rect 9823 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10139 8736
rect 9823 8671 10139 8672
rect 14262 8736 14578 8737
rect 14262 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14578 8736
rect 14262 8671 14578 8672
rect 18701 8736 19017 8737
rect 18701 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19017 8736
rect 19200 8712 20000 8742
rect 18701 8671 19017 8672
rect 0 8440 800 8560
rect 16246 8468 16252 8532
rect 16316 8530 16322 8532
rect 17033 8530 17099 8533
rect 16316 8528 17099 8530
rect 16316 8472 17038 8528
rect 17094 8472 17099 8528
rect 16316 8470 17099 8472
rect 16316 8468 16322 8470
rect 17033 8467 17099 8470
rect 19200 8304 20000 8424
rect 3165 8192 3481 8193
rect 0 8122 800 8152
rect 3165 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3481 8192
rect 3165 8127 3481 8128
rect 7604 8192 7920 8193
rect 7604 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7920 8192
rect 7604 8127 7920 8128
rect 12043 8192 12359 8193
rect 12043 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12359 8192
rect 12043 8127 12359 8128
rect 16482 8192 16798 8193
rect 16482 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16798 8192
rect 16482 8127 16798 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 800 8062
rect 1577 8059 1643 8062
rect 18321 7986 18387 7989
rect 19200 7986 20000 8016
rect 18321 7984 20000 7986
rect 18321 7928 18326 7984
rect 18382 7928 20000 7984
rect 18321 7926 20000 7928
rect 18321 7923 18387 7926
rect 19200 7896 20000 7926
rect 0 7714 800 7744
rect 1577 7714 1643 7717
rect 0 7712 1643 7714
rect 0 7656 1582 7712
rect 1638 7656 1643 7712
rect 0 7654 1643 7656
rect 0 7624 800 7654
rect 1577 7651 1643 7654
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 19200 7578 20000 7608
rect 19152 7488 20000 7578
rect 18321 7442 18387 7445
rect 19152 7442 19212 7488
rect 18321 7440 19212 7442
rect 18321 7384 18326 7440
rect 18382 7384 19212 7440
rect 18321 7382 19212 7384
rect 18321 7379 18387 7382
rect 0 7216 800 7336
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 19200 7080 20000 7200
rect 16482 7039 16798 7040
rect 0 6898 800 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 800 6838
rect 1577 6835 1643 6838
rect 18321 6762 18387 6765
rect 19200 6762 20000 6792
rect 18321 6760 20000 6762
rect 18321 6704 18326 6760
rect 18382 6704 20000 6760
rect 18321 6702 20000 6704
rect 18321 6699 18387 6702
rect 19200 6672 20000 6702
rect 5384 6560 5700 6561
rect 0 6490 800 6520
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 1577 6490 1643 6493
rect 0 6488 1643 6490
rect 0 6432 1582 6488
rect 1638 6432 1643 6488
rect 0 6430 1643 6432
rect 0 6400 800 6430
rect 1577 6427 1643 6430
rect 18321 6354 18387 6357
rect 19200 6354 20000 6384
rect 18321 6352 20000 6354
rect 18321 6296 18326 6352
rect 18382 6296 20000 6352
rect 18321 6294 20000 6296
rect 18321 6291 18387 6294
rect 19200 6264 20000 6294
rect 0 5992 800 6112
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 19200 5856 20000 5976
rect 0 5674 800 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 800 5614
rect 1577 5611 1643 5614
rect 18321 5674 18387 5677
rect 18321 5672 19212 5674
rect 18321 5616 18326 5672
rect 18382 5616 19212 5672
rect 18321 5614 19212 5616
rect 18321 5611 18387 5614
rect 19152 5568 19212 5614
rect 19152 5478 20000 5568
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 19200 5448 20000 5478
rect 18701 5407 19017 5408
rect 0 5266 800 5296
rect 1577 5266 1643 5269
rect 0 5264 1643 5266
rect 0 5208 1582 5264
rect 1638 5208 1643 5264
rect 0 5206 1643 5208
rect 0 5176 800 5206
rect 1577 5203 1643 5206
rect 18321 5130 18387 5133
rect 19200 5130 20000 5160
rect 18321 5128 20000 5130
rect 18321 5072 18326 5128
rect 18382 5072 20000 5128
rect 18321 5070 20000 5072
rect 18321 5067 18387 5070
rect 19200 5040 20000 5070
rect 3165 4928 3481 4929
rect 0 4768 800 4888
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 19200 4632 20000 4752
rect 0 4450 800 4480
rect 1577 4450 1643 4453
rect 0 4448 1643 4450
rect 0 4392 1582 4448
rect 1638 4392 1643 4448
rect 0 4390 1643 4392
rect 0 4360 800 4390
rect 1577 4387 1643 4390
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 19200 4317 20000 4344
rect 19149 4312 20000 4317
rect 19149 4256 19154 4312
rect 19210 4256 20000 4312
rect 19149 4251 20000 4256
rect 19200 4224 20000 4251
rect 0 4042 800 4072
rect 1577 4042 1643 4045
rect 0 4040 1643 4042
rect 0 3984 1582 4040
rect 1638 3984 1643 4040
rect 0 3982 1643 3984
rect 0 3952 800 3982
rect 1577 3979 1643 3982
rect 18321 3906 18387 3909
rect 19200 3906 20000 3936
rect 18321 3904 20000 3906
rect 18321 3848 18326 3904
rect 18382 3848 20000 3904
rect 18321 3846 20000 3848
rect 18321 3843 18387 3846
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 19200 3816 20000 3846
rect 16482 3775 16798 3776
rect 0 3544 800 3664
rect 19200 3408 20000 3528
rect 5384 3296 5700 3297
rect 0 3226 800 3256
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 1577 3226 1643 3229
rect 0 3224 1643 3226
rect 0 3168 1582 3224
rect 1638 3168 1643 3224
rect 0 3166 1643 3168
rect 0 3136 800 3166
rect 1577 3163 1643 3166
rect 18321 3090 18387 3093
rect 19200 3090 20000 3120
rect 18321 3088 20000 3090
rect 18321 3032 18326 3088
rect 18382 3032 20000 3088
rect 18321 3030 20000 3032
rect 18321 3027 18387 3030
rect 19200 3000 20000 3030
rect 0 2818 800 2848
rect 1577 2818 1643 2821
rect 0 2816 1643 2818
rect 0 2760 1582 2816
rect 1638 2760 1643 2816
rect 0 2758 1643 2760
rect 0 2728 800 2758
rect 1577 2755 1643 2758
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 18321 2682 18387 2685
rect 19200 2682 20000 2712
rect 18321 2680 20000 2682
rect 18321 2624 18326 2680
rect 18382 2624 20000 2680
rect 18321 2622 20000 2624
rect 18321 2619 18387 2622
rect 19200 2592 20000 2622
rect 0 2320 800 2440
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 19200 2184 20000 2304
rect 18701 2143 19017 2144
rect 0 2002 800 2032
rect 2221 2002 2287 2005
rect 0 2000 2287 2002
rect 0 1944 2226 2000
rect 2282 1944 2287 2000
rect 0 1942 2287 1944
rect 0 1912 800 1942
rect 2221 1939 2287 1942
rect 18321 1866 18387 1869
rect 19200 1866 20000 1896
rect 18321 1864 20000 1866
rect 18321 1808 18326 1864
rect 18382 1808 20000 1864
rect 18321 1806 20000 1808
rect 18321 1803 18387 1806
rect 19200 1776 20000 1806
rect 0 1594 800 1624
rect 1577 1594 1643 1597
rect 0 1592 1643 1594
rect 0 1536 1582 1592
rect 1638 1536 1643 1592
rect 0 1534 1643 1536
rect 0 1504 800 1534
rect 1577 1531 1643 1534
rect 17677 1458 17743 1461
rect 19200 1458 20000 1488
rect 17677 1456 20000 1458
rect 17677 1400 17682 1456
rect 17738 1400 20000 1456
rect 17677 1398 20000 1400
rect 17677 1395 17743 1398
rect 19200 1368 20000 1398
rect 19200 960 20000 1080
<< via3 >>
rect 16252 18532 16316 18596
rect 5390 17436 5454 17440
rect 5390 17380 5394 17436
rect 5394 17380 5450 17436
rect 5450 17380 5454 17436
rect 5390 17376 5454 17380
rect 5470 17436 5534 17440
rect 5470 17380 5474 17436
rect 5474 17380 5530 17436
rect 5530 17380 5534 17436
rect 5470 17376 5534 17380
rect 5550 17436 5614 17440
rect 5550 17380 5554 17436
rect 5554 17380 5610 17436
rect 5610 17380 5614 17436
rect 5550 17376 5614 17380
rect 5630 17436 5694 17440
rect 5630 17380 5634 17436
rect 5634 17380 5690 17436
rect 5690 17380 5694 17436
rect 5630 17376 5694 17380
rect 9829 17436 9893 17440
rect 9829 17380 9833 17436
rect 9833 17380 9889 17436
rect 9889 17380 9893 17436
rect 9829 17376 9893 17380
rect 9909 17436 9973 17440
rect 9909 17380 9913 17436
rect 9913 17380 9969 17436
rect 9969 17380 9973 17436
rect 9909 17376 9973 17380
rect 9989 17436 10053 17440
rect 9989 17380 9993 17436
rect 9993 17380 10049 17436
rect 10049 17380 10053 17436
rect 9989 17376 10053 17380
rect 10069 17436 10133 17440
rect 10069 17380 10073 17436
rect 10073 17380 10129 17436
rect 10129 17380 10133 17436
rect 10069 17376 10133 17380
rect 14268 17436 14332 17440
rect 14268 17380 14272 17436
rect 14272 17380 14328 17436
rect 14328 17380 14332 17436
rect 14268 17376 14332 17380
rect 14348 17436 14412 17440
rect 14348 17380 14352 17436
rect 14352 17380 14408 17436
rect 14408 17380 14412 17436
rect 14348 17376 14412 17380
rect 14428 17436 14492 17440
rect 14428 17380 14432 17436
rect 14432 17380 14488 17436
rect 14488 17380 14492 17436
rect 14428 17376 14492 17380
rect 14508 17436 14572 17440
rect 14508 17380 14512 17436
rect 14512 17380 14568 17436
rect 14568 17380 14572 17436
rect 14508 17376 14572 17380
rect 18707 17436 18771 17440
rect 18707 17380 18711 17436
rect 18711 17380 18767 17436
rect 18767 17380 18771 17436
rect 18707 17376 18771 17380
rect 18787 17436 18851 17440
rect 18787 17380 18791 17436
rect 18791 17380 18847 17436
rect 18847 17380 18851 17436
rect 18787 17376 18851 17380
rect 18867 17436 18931 17440
rect 18867 17380 18871 17436
rect 18871 17380 18927 17436
rect 18927 17380 18931 17436
rect 18867 17376 18931 17380
rect 18947 17436 19011 17440
rect 18947 17380 18951 17436
rect 18951 17380 19007 17436
rect 19007 17380 19011 17436
rect 18947 17376 19011 17380
rect 3171 16892 3235 16896
rect 3171 16836 3175 16892
rect 3175 16836 3231 16892
rect 3231 16836 3235 16892
rect 3171 16832 3235 16836
rect 3251 16892 3315 16896
rect 3251 16836 3255 16892
rect 3255 16836 3311 16892
rect 3311 16836 3315 16892
rect 3251 16832 3315 16836
rect 3331 16892 3395 16896
rect 3331 16836 3335 16892
rect 3335 16836 3391 16892
rect 3391 16836 3395 16892
rect 3331 16832 3395 16836
rect 3411 16892 3475 16896
rect 3411 16836 3415 16892
rect 3415 16836 3471 16892
rect 3471 16836 3475 16892
rect 3411 16832 3475 16836
rect 7610 16892 7674 16896
rect 7610 16836 7614 16892
rect 7614 16836 7670 16892
rect 7670 16836 7674 16892
rect 7610 16832 7674 16836
rect 7690 16892 7754 16896
rect 7690 16836 7694 16892
rect 7694 16836 7750 16892
rect 7750 16836 7754 16892
rect 7690 16832 7754 16836
rect 7770 16892 7834 16896
rect 7770 16836 7774 16892
rect 7774 16836 7830 16892
rect 7830 16836 7834 16892
rect 7770 16832 7834 16836
rect 7850 16892 7914 16896
rect 7850 16836 7854 16892
rect 7854 16836 7910 16892
rect 7910 16836 7914 16892
rect 7850 16832 7914 16836
rect 12049 16892 12113 16896
rect 12049 16836 12053 16892
rect 12053 16836 12109 16892
rect 12109 16836 12113 16892
rect 12049 16832 12113 16836
rect 12129 16892 12193 16896
rect 12129 16836 12133 16892
rect 12133 16836 12189 16892
rect 12189 16836 12193 16892
rect 12129 16832 12193 16836
rect 12209 16892 12273 16896
rect 12209 16836 12213 16892
rect 12213 16836 12269 16892
rect 12269 16836 12273 16892
rect 12209 16832 12273 16836
rect 12289 16892 12353 16896
rect 12289 16836 12293 16892
rect 12293 16836 12349 16892
rect 12349 16836 12353 16892
rect 12289 16832 12353 16836
rect 16488 16892 16552 16896
rect 16488 16836 16492 16892
rect 16492 16836 16548 16892
rect 16548 16836 16552 16892
rect 16488 16832 16552 16836
rect 16568 16892 16632 16896
rect 16568 16836 16572 16892
rect 16572 16836 16628 16892
rect 16628 16836 16632 16892
rect 16568 16832 16632 16836
rect 16648 16892 16712 16896
rect 16648 16836 16652 16892
rect 16652 16836 16708 16892
rect 16708 16836 16712 16892
rect 16648 16832 16712 16836
rect 16728 16892 16792 16896
rect 16728 16836 16732 16892
rect 16732 16836 16788 16892
rect 16788 16836 16792 16892
rect 16728 16832 16792 16836
rect 5390 16348 5454 16352
rect 5390 16292 5394 16348
rect 5394 16292 5450 16348
rect 5450 16292 5454 16348
rect 5390 16288 5454 16292
rect 5470 16348 5534 16352
rect 5470 16292 5474 16348
rect 5474 16292 5530 16348
rect 5530 16292 5534 16348
rect 5470 16288 5534 16292
rect 5550 16348 5614 16352
rect 5550 16292 5554 16348
rect 5554 16292 5610 16348
rect 5610 16292 5614 16348
rect 5550 16288 5614 16292
rect 5630 16348 5694 16352
rect 5630 16292 5634 16348
rect 5634 16292 5690 16348
rect 5690 16292 5694 16348
rect 5630 16288 5694 16292
rect 9829 16348 9893 16352
rect 9829 16292 9833 16348
rect 9833 16292 9889 16348
rect 9889 16292 9893 16348
rect 9829 16288 9893 16292
rect 9909 16348 9973 16352
rect 9909 16292 9913 16348
rect 9913 16292 9969 16348
rect 9969 16292 9973 16348
rect 9909 16288 9973 16292
rect 9989 16348 10053 16352
rect 9989 16292 9993 16348
rect 9993 16292 10049 16348
rect 10049 16292 10053 16348
rect 9989 16288 10053 16292
rect 10069 16348 10133 16352
rect 10069 16292 10073 16348
rect 10073 16292 10129 16348
rect 10129 16292 10133 16348
rect 10069 16288 10133 16292
rect 14268 16348 14332 16352
rect 14268 16292 14272 16348
rect 14272 16292 14328 16348
rect 14328 16292 14332 16348
rect 14268 16288 14332 16292
rect 14348 16348 14412 16352
rect 14348 16292 14352 16348
rect 14352 16292 14408 16348
rect 14408 16292 14412 16348
rect 14348 16288 14412 16292
rect 14428 16348 14492 16352
rect 14428 16292 14432 16348
rect 14432 16292 14488 16348
rect 14488 16292 14492 16348
rect 14428 16288 14492 16292
rect 14508 16348 14572 16352
rect 14508 16292 14512 16348
rect 14512 16292 14568 16348
rect 14568 16292 14572 16348
rect 14508 16288 14572 16292
rect 15884 16280 15948 16284
rect 15884 16224 15898 16280
rect 15898 16224 15948 16280
rect 15884 16220 15948 16224
rect 10548 16084 10612 16148
rect 18707 16348 18771 16352
rect 18707 16292 18711 16348
rect 18711 16292 18767 16348
rect 18767 16292 18771 16348
rect 18707 16288 18771 16292
rect 18787 16348 18851 16352
rect 18787 16292 18791 16348
rect 18791 16292 18847 16348
rect 18847 16292 18851 16348
rect 18787 16288 18851 16292
rect 18867 16348 18931 16352
rect 18867 16292 18871 16348
rect 18871 16292 18927 16348
rect 18927 16292 18931 16348
rect 18867 16288 18931 16292
rect 18947 16348 19011 16352
rect 18947 16292 18951 16348
rect 18951 16292 19007 16348
rect 19007 16292 19011 16348
rect 18947 16288 19011 16292
rect 3171 15804 3235 15808
rect 3171 15748 3175 15804
rect 3175 15748 3231 15804
rect 3231 15748 3235 15804
rect 3171 15744 3235 15748
rect 3251 15804 3315 15808
rect 3251 15748 3255 15804
rect 3255 15748 3311 15804
rect 3311 15748 3315 15804
rect 3251 15744 3315 15748
rect 3331 15804 3395 15808
rect 3331 15748 3335 15804
rect 3335 15748 3391 15804
rect 3391 15748 3395 15804
rect 3331 15744 3395 15748
rect 3411 15804 3475 15808
rect 3411 15748 3415 15804
rect 3415 15748 3471 15804
rect 3471 15748 3475 15804
rect 3411 15744 3475 15748
rect 7610 15804 7674 15808
rect 7610 15748 7614 15804
rect 7614 15748 7670 15804
rect 7670 15748 7674 15804
rect 7610 15744 7674 15748
rect 7690 15804 7754 15808
rect 7690 15748 7694 15804
rect 7694 15748 7750 15804
rect 7750 15748 7754 15804
rect 7690 15744 7754 15748
rect 7770 15804 7834 15808
rect 7770 15748 7774 15804
rect 7774 15748 7830 15804
rect 7830 15748 7834 15804
rect 7770 15744 7834 15748
rect 7850 15804 7914 15808
rect 7850 15748 7854 15804
rect 7854 15748 7910 15804
rect 7910 15748 7914 15804
rect 7850 15744 7914 15748
rect 12049 15804 12113 15808
rect 12049 15748 12053 15804
rect 12053 15748 12109 15804
rect 12109 15748 12113 15804
rect 12049 15744 12113 15748
rect 12129 15804 12193 15808
rect 12129 15748 12133 15804
rect 12133 15748 12189 15804
rect 12189 15748 12193 15804
rect 12129 15744 12193 15748
rect 12209 15804 12273 15808
rect 12209 15748 12213 15804
rect 12213 15748 12269 15804
rect 12269 15748 12273 15804
rect 12209 15744 12273 15748
rect 12289 15804 12353 15808
rect 12289 15748 12293 15804
rect 12293 15748 12349 15804
rect 12349 15748 12353 15804
rect 12289 15744 12353 15748
rect 16488 15804 16552 15808
rect 16488 15748 16492 15804
rect 16492 15748 16548 15804
rect 16548 15748 16552 15804
rect 16488 15744 16552 15748
rect 16568 15804 16632 15808
rect 16568 15748 16572 15804
rect 16572 15748 16628 15804
rect 16628 15748 16632 15804
rect 16568 15744 16632 15748
rect 16648 15804 16712 15808
rect 16648 15748 16652 15804
rect 16652 15748 16708 15804
rect 16708 15748 16712 15804
rect 16648 15744 16712 15748
rect 16728 15804 16792 15808
rect 16728 15748 16732 15804
rect 16732 15748 16788 15804
rect 16788 15748 16792 15804
rect 16728 15744 16792 15748
rect 11100 15540 11164 15604
rect 13860 15540 13924 15604
rect 5390 15260 5454 15264
rect 5390 15204 5394 15260
rect 5394 15204 5450 15260
rect 5450 15204 5454 15260
rect 5390 15200 5454 15204
rect 5470 15260 5534 15264
rect 5470 15204 5474 15260
rect 5474 15204 5530 15260
rect 5530 15204 5534 15260
rect 5470 15200 5534 15204
rect 5550 15260 5614 15264
rect 5550 15204 5554 15260
rect 5554 15204 5610 15260
rect 5610 15204 5614 15260
rect 5550 15200 5614 15204
rect 5630 15260 5694 15264
rect 5630 15204 5634 15260
rect 5634 15204 5690 15260
rect 5690 15204 5694 15260
rect 5630 15200 5694 15204
rect 9829 15260 9893 15264
rect 9829 15204 9833 15260
rect 9833 15204 9889 15260
rect 9889 15204 9893 15260
rect 9829 15200 9893 15204
rect 9909 15260 9973 15264
rect 9909 15204 9913 15260
rect 9913 15204 9969 15260
rect 9969 15204 9973 15260
rect 9909 15200 9973 15204
rect 9989 15260 10053 15264
rect 9989 15204 9993 15260
rect 9993 15204 10049 15260
rect 10049 15204 10053 15260
rect 9989 15200 10053 15204
rect 10069 15260 10133 15264
rect 10069 15204 10073 15260
rect 10073 15204 10129 15260
rect 10129 15204 10133 15260
rect 10069 15200 10133 15204
rect 14268 15260 14332 15264
rect 14268 15204 14272 15260
rect 14272 15204 14328 15260
rect 14328 15204 14332 15260
rect 14268 15200 14332 15204
rect 14348 15260 14412 15264
rect 14348 15204 14352 15260
rect 14352 15204 14408 15260
rect 14408 15204 14412 15260
rect 14348 15200 14412 15204
rect 14428 15260 14492 15264
rect 14428 15204 14432 15260
rect 14432 15204 14488 15260
rect 14488 15204 14492 15260
rect 14428 15200 14492 15204
rect 14508 15260 14572 15264
rect 14508 15204 14512 15260
rect 14512 15204 14568 15260
rect 14568 15204 14572 15260
rect 14508 15200 14572 15204
rect 18707 15260 18771 15264
rect 18707 15204 18711 15260
rect 18711 15204 18767 15260
rect 18767 15204 18771 15260
rect 18707 15200 18771 15204
rect 18787 15260 18851 15264
rect 18787 15204 18791 15260
rect 18791 15204 18847 15260
rect 18847 15204 18851 15260
rect 18787 15200 18851 15204
rect 18867 15260 18931 15264
rect 18867 15204 18871 15260
rect 18871 15204 18927 15260
rect 18927 15204 18931 15260
rect 18867 15200 18931 15204
rect 18947 15260 19011 15264
rect 18947 15204 18951 15260
rect 18951 15204 19007 15260
rect 19007 15204 19011 15260
rect 18947 15200 19011 15204
rect 3171 14716 3235 14720
rect 3171 14660 3175 14716
rect 3175 14660 3231 14716
rect 3231 14660 3235 14716
rect 3171 14656 3235 14660
rect 3251 14716 3315 14720
rect 3251 14660 3255 14716
rect 3255 14660 3311 14716
rect 3311 14660 3315 14716
rect 3251 14656 3315 14660
rect 3331 14716 3395 14720
rect 3331 14660 3335 14716
rect 3335 14660 3391 14716
rect 3391 14660 3395 14716
rect 3331 14656 3395 14660
rect 3411 14716 3475 14720
rect 3411 14660 3415 14716
rect 3415 14660 3471 14716
rect 3471 14660 3475 14716
rect 3411 14656 3475 14660
rect 7610 14716 7674 14720
rect 7610 14660 7614 14716
rect 7614 14660 7670 14716
rect 7670 14660 7674 14716
rect 7610 14656 7674 14660
rect 7690 14716 7754 14720
rect 7690 14660 7694 14716
rect 7694 14660 7750 14716
rect 7750 14660 7754 14716
rect 7690 14656 7754 14660
rect 7770 14716 7834 14720
rect 7770 14660 7774 14716
rect 7774 14660 7830 14716
rect 7830 14660 7834 14716
rect 7770 14656 7834 14660
rect 7850 14716 7914 14720
rect 7850 14660 7854 14716
rect 7854 14660 7910 14716
rect 7910 14660 7914 14716
rect 7850 14656 7914 14660
rect 12049 14716 12113 14720
rect 12049 14660 12053 14716
rect 12053 14660 12109 14716
rect 12109 14660 12113 14716
rect 12049 14656 12113 14660
rect 12129 14716 12193 14720
rect 12129 14660 12133 14716
rect 12133 14660 12189 14716
rect 12189 14660 12193 14716
rect 12129 14656 12193 14660
rect 12209 14716 12273 14720
rect 12209 14660 12213 14716
rect 12213 14660 12269 14716
rect 12269 14660 12273 14716
rect 12209 14656 12273 14660
rect 12289 14716 12353 14720
rect 12289 14660 12293 14716
rect 12293 14660 12349 14716
rect 12349 14660 12353 14716
rect 12289 14656 12353 14660
rect 16488 14716 16552 14720
rect 16488 14660 16492 14716
rect 16492 14660 16548 14716
rect 16548 14660 16552 14716
rect 16488 14656 16552 14660
rect 16568 14716 16632 14720
rect 16568 14660 16572 14716
rect 16572 14660 16628 14716
rect 16628 14660 16632 14716
rect 16568 14656 16632 14660
rect 16648 14716 16712 14720
rect 16648 14660 16652 14716
rect 16652 14660 16708 14716
rect 16708 14660 16712 14716
rect 16648 14656 16712 14660
rect 16728 14716 16792 14720
rect 16728 14660 16732 14716
rect 16732 14660 16788 14716
rect 16788 14660 16792 14716
rect 16728 14656 16792 14660
rect 12940 14452 13004 14516
rect 16068 14452 16132 14516
rect 5390 14172 5454 14176
rect 5390 14116 5394 14172
rect 5394 14116 5450 14172
rect 5450 14116 5454 14172
rect 5390 14112 5454 14116
rect 5470 14172 5534 14176
rect 5470 14116 5474 14172
rect 5474 14116 5530 14172
rect 5530 14116 5534 14172
rect 5470 14112 5534 14116
rect 5550 14172 5614 14176
rect 5550 14116 5554 14172
rect 5554 14116 5610 14172
rect 5610 14116 5614 14172
rect 5550 14112 5614 14116
rect 5630 14172 5694 14176
rect 5630 14116 5634 14172
rect 5634 14116 5690 14172
rect 5690 14116 5694 14172
rect 5630 14112 5694 14116
rect 9829 14172 9893 14176
rect 9829 14116 9833 14172
rect 9833 14116 9889 14172
rect 9889 14116 9893 14172
rect 9829 14112 9893 14116
rect 9909 14172 9973 14176
rect 9909 14116 9913 14172
rect 9913 14116 9969 14172
rect 9969 14116 9973 14172
rect 9909 14112 9973 14116
rect 9989 14172 10053 14176
rect 9989 14116 9993 14172
rect 9993 14116 10049 14172
rect 10049 14116 10053 14172
rect 9989 14112 10053 14116
rect 10069 14172 10133 14176
rect 10069 14116 10073 14172
rect 10073 14116 10129 14172
rect 10129 14116 10133 14172
rect 10069 14112 10133 14116
rect 14268 14172 14332 14176
rect 14268 14116 14272 14172
rect 14272 14116 14328 14172
rect 14328 14116 14332 14172
rect 14268 14112 14332 14116
rect 14348 14172 14412 14176
rect 14348 14116 14352 14172
rect 14352 14116 14408 14172
rect 14408 14116 14412 14172
rect 14348 14112 14412 14116
rect 14428 14172 14492 14176
rect 14428 14116 14432 14172
rect 14432 14116 14488 14172
rect 14488 14116 14492 14172
rect 14428 14112 14492 14116
rect 14508 14172 14572 14176
rect 14508 14116 14512 14172
rect 14512 14116 14568 14172
rect 14568 14116 14572 14172
rect 14508 14112 14572 14116
rect 18707 14172 18771 14176
rect 18707 14116 18711 14172
rect 18711 14116 18767 14172
rect 18767 14116 18771 14172
rect 18707 14112 18771 14116
rect 18787 14172 18851 14176
rect 18787 14116 18791 14172
rect 18791 14116 18847 14172
rect 18847 14116 18851 14172
rect 18787 14112 18851 14116
rect 18867 14172 18931 14176
rect 18867 14116 18871 14172
rect 18871 14116 18927 14172
rect 18927 14116 18931 14172
rect 18867 14112 18931 14116
rect 18947 14172 19011 14176
rect 18947 14116 18951 14172
rect 18951 14116 19007 14172
rect 19007 14116 19011 14172
rect 18947 14112 19011 14116
rect 11100 14044 11164 14108
rect 15700 13772 15764 13836
rect 12940 13696 13004 13700
rect 12940 13640 12954 13696
rect 12954 13640 13004 13696
rect 12940 13636 13004 13640
rect 3171 13628 3235 13632
rect 3171 13572 3175 13628
rect 3175 13572 3231 13628
rect 3231 13572 3235 13628
rect 3171 13568 3235 13572
rect 3251 13628 3315 13632
rect 3251 13572 3255 13628
rect 3255 13572 3311 13628
rect 3311 13572 3315 13628
rect 3251 13568 3315 13572
rect 3331 13628 3395 13632
rect 3331 13572 3335 13628
rect 3335 13572 3391 13628
rect 3391 13572 3395 13628
rect 3331 13568 3395 13572
rect 3411 13628 3475 13632
rect 3411 13572 3415 13628
rect 3415 13572 3471 13628
rect 3471 13572 3475 13628
rect 3411 13568 3475 13572
rect 7610 13628 7674 13632
rect 7610 13572 7614 13628
rect 7614 13572 7670 13628
rect 7670 13572 7674 13628
rect 7610 13568 7674 13572
rect 7690 13628 7754 13632
rect 7690 13572 7694 13628
rect 7694 13572 7750 13628
rect 7750 13572 7754 13628
rect 7690 13568 7754 13572
rect 7770 13628 7834 13632
rect 7770 13572 7774 13628
rect 7774 13572 7830 13628
rect 7830 13572 7834 13628
rect 7770 13568 7834 13572
rect 7850 13628 7914 13632
rect 7850 13572 7854 13628
rect 7854 13572 7910 13628
rect 7910 13572 7914 13628
rect 7850 13568 7914 13572
rect 12049 13628 12113 13632
rect 12049 13572 12053 13628
rect 12053 13572 12109 13628
rect 12109 13572 12113 13628
rect 12049 13568 12113 13572
rect 12129 13628 12193 13632
rect 12129 13572 12133 13628
rect 12133 13572 12189 13628
rect 12189 13572 12193 13628
rect 12129 13568 12193 13572
rect 12209 13628 12273 13632
rect 12209 13572 12213 13628
rect 12213 13572 12269 13628
rect 12269 13572 12273 13628
rect 12209 13568 12273 13572
rect 12289 13628 12353 13632
rect 12289 13572 12293 13628
rect 12293 13572 12349 13628
rect 12349 13572 12353 13628
rect 12289 13568 12353 13572
rect 16488 13628 16552 13632
rect 16488 13572 16492 13628
rect 16492 13572 16548 13628
rect 16548 13572 16552 13628
rect 16488 13568 16552 13572
rect 16568 13628 16632 13632
rect 16568 13572 16572 13628
rect 16572 13572 16628 13628
rect 16628 13572 16632 13628
rect 16568 13568 16632 13572
rect 16648 13628 16712 13632
rect 16648 13572 16652 13628
rect 16652 13572 16708 13628
rect 16708 13572 16712 13628
rect 16648 13568 16712 13572
rect 16728 13628 16792 13632
rect 16728 13572 16732 13628
rect 16732 13572 16788 13628
rect 16788 13572 16792 13628
rect 16728 13568 16792 13572
rect 16988 13288 17052 13292
rect 16988 13232 17038 13288
rect 17038 13232 17052 13288
rect 16988 13228 17052 13232
rect 5390 13084 5454 13088
rect 5390 13028 5394 13084
rect 5394 13028 5450 13084
rect 5450 13028 5454 13084
rect 5390 13024 5454 13028
rect 5470 13084 5534 13088
rect 5470 13028 5474 13084
rect 5474 13028 5530 13084
rect 5530 13028 5534 13084
rect 5470 13024 5534 13028
rect 5550 13084 5614 13088
rect 5550 13028 5554 13084
rect 5554 13028 5610 13084
rect 5610 13028 5614 13084
rect 5550 13024 5614 13028
rect 5630 13084 5694 13088
rect 5630 13028 5634 13084
rect 5634 13028 5690 13084
rect 5690 13028 5694 13084
rect 5630 13024 5694 13028
rect 9829 13084 9893 13088
rect 9829 13028 9833 13084
rect 9833 13028 9889 13084
rect 9889 13028 9893 13084
rect 9829 13024 9893 13028
rect 9909 13084 9973 13088
rect 9909 13028 9913 13084
rect 9913 13028 9969 13084
rect 9969 13028 9973 13084
rect 9909 13024 9973 13028
rect 9989 13084 10053 13088
rect 9989 13028 9993 13084
rect 9993 13028 10049 13084
rect 10049 13028 10053 13084
rect 9989 13024 10053 13028
rect 10069 13084 10133 13088
rect 10069 13028 10073 13084
rect 10073 13028 10129 13084
rect 10129 13028 10133 13084
rect 10069 13024 10133 13028
rect 14268 13084 14332 13088
rect 14268 13028 14272 13084
rect 14272 13028 14328 13084
rect 14328 13028 14332 13084
rect 14268 13024 14332 13028
rect 14348 13084 14412 13088
rect 14348 13028 14352 13084
rect 14352 13028 14408 13084
rect 14408 13028 14412 13084
rect 14348 13024 14412 13028
rect 14428 13084 14492 13088
rect 14428 13028 14432 13084
rect 14432 13028 14488 13084
rect 14488 13028 14492 13084
rect 14428 13024 14492 13028
rect 14508 13084 14572 13088
rect 14508 13028 14512 13084
rect 14512 13028 14568 13084
rect 14568 13028 14572 13084
rect 14508 13024 14572 13028
rect 18707 13084 18771 13088
rect 18707 13028 18711 13084
rect 18711 13028 18767 13084
rect 18767 13028 18771 13084
rect 18707 13024 18771 13028
rect 18787 13084 18851 13088
rect 18787 13028 18791 13084
rect 18791 13028 18847 13084
rect 18847 13028 18851 13084
rect 18787 13024 18851 13028
rect 18867 13084 18931 13088
rect 18867 13028 18871 13084
rect 18871 13028 18927 13084
rect 18927 13028 18931 13084
rect 18867 13024 18931 13028
rect 18947 13084 19011 13088
rect 18947 13028 18951 13084
rect 18951 13028 19007 13084
rect 19007 13028 19011 13084
rect 18947 13024 19011 13028
rect 10548 12880 10612 12884
rect 10548 12824 10562 12880
rect 10562 12824 10612 12880
rect 10548 12820 10612 12824
rect 3171 12540 3235 12544
rect 3171 12484 3175 12540
rect 3175 12484 3231 12540
rect 3231 12484 3235 12540
rect 3171 12480 3235 12484
rect 3251 12540 3315 12544
rect 3251 12484 3255 12540
rect 3255 12484 3311 12540
rect 3311 12484 3315 12540
rect 3251 12480 3315 12484
rect 3331 12540 3395 12544
rect 3331 12484 3335 12540
rect 3335 12484 3391 12540
rect 3391 12484 3395 12540
rect 3331 12480 3395 12484
rect 3411 12540 3475 12544
rect 3411 12484 3415 12540
rect 3415 12484 3471 12540
rect 3471 12484 3475 12540
rect 3411 12480 3475 12484
rect 7610 12540 7674 12544
rect 7610 12484 7614 12540
rect 7614 12484 7670 12540
rect 7670 12484 7674 12540
rect 7610 12480 7674 12484
rect 7690 12540 7754 12544
rect 7690 12484 7694 12540
rect 7694 12484 7750 12540
rect 7750 12484 7754 12540
rect 7690 12480 7754 12484
rect 7770 12540 7834 12544
rect 7770 12484 7774 12540
rect 7774 12484 7830 12540
rect 7830 12484 7834 12540
rect 7770 12480 7834 12484
rect 7850 12540 7914 12544
rect 7850 12484 7854 12540
rect 7854 12484 7910 12540
rect 7910 12484 7914 12540
rect 7850 12480 7914 12484
rect 12049 12540 12113 12544
rect 12049 12484 12053 12540
rect 12053 12484 12109 12540
rect 12109 12484 12113 12540
rect 12049 12480 12113 12484
rect 12129 12540 12193 12544
rect 12129 12484 12133 12540
rect 12133 12484 12189 12540
rect 12189 12484 12193 12540
rect 12129 12480 12193 12484
rect 12209 12540 12273 12544
rect 12209 12484 12213 12540
rect 12213 12484 12269 12540
rect 12269 12484 12273 12540
rect 12209 12480 12273 12484
rect 12289 12540 12353 12544
rect 12289 12484 12293 12540
rect 12293 12484 12349 12540
rect 12349 12484 12353 12540
rect 12289 12480 12353 12484
rect 16488 12540 16552 12544
rect 16488 12484 16492 12540
rect 16492 12484 16548 12540
rect 16548 12484 16552 12540
rect 16488 12480 16552 12484
rect 16568 12540 16632 12544
rect 16568 12484 16572 12540
rect 16572 12484 16628 12540
rect 16628 12484 16632 12540
rect 16568 12480 16632 12484
rect 16648 12540 16712 12544
rect 16648 12484 16652 12540
rect 16652 12484 16708 12540
rect 16708 12484 16712 12540
rect 16648 12480 16712 12484
rect 16728 12540 16792 12544
rect 16728 12484 16732 12540
rect 16732 12484 16788 12540
rect 16788 12484 16792 12540
rect 16728 12480 16792 12484
rect 16068 12472 16132 12476
rect 16068 12416 16118 12472
rect 16118 12416 16132 12472
rect 16068 12412 16132 12416
rect 15884 12004 15948 12068
rect 5390 11996 5454 12000
rect 5390 11940 5394 11996
rect 5394 11940 5450 11996
rect 5450 11940 5454 11996
rect 5390 11936 5454 11940
rect 5470 11996 5534 12000
rect 5470 11940 5474 11996
rect 5474 11940 5530 11996
rect 5530 11940 5534 11996
rect 5470 11936 5534 11940
rect 5550 11996 5614 12000
rect 5550 11940 5554 11996
rect 5554 11940 5610 11996
rect 5610 11940 5614 11996
rect 5550 11936 5614 11940
rect 5630 11996 5694 12000
rect 5630 11940 5634 11996
rect 5634 11940 5690 11996
rect 5690 11940 5694 11996
rect 5630 11936 5694 11940
rect 9829 11996 9893 12000
rect 9829 11940 9833 11996
rect 9833 11940 9889 11996
rect 9889 11940 9893 11996
rect 9829 11936 9893 11940
rect 9909 11996 9973 12000
rect 9909 11940 9913 11996
rect 9913 11940 9969 11996
rect 9969 11940 9973 11996
rect 9909 11936 9973 11940
rect 9989 11996 10053 12000
rect 9989 11940 9993 11996
rect 9993 11940 10049 11996
rect 10049 11940 10053 11996
rect 9989 11936 10053 11940
rect 10069 11996 10133 12000
rect 10069 11940 10073 11996
rect 10073 11940 10129 11996
rect 10129 11940 10133 11996
rect 10069 11936 10133 11940
rect 14268 11996 14332 12000
rect 14268 11940 14272 11996
rect 14272 11940 14328 11996
rect 14328 11940 14332 11996
rect 14268 11936 14332 11940
rect 14348 11996 14412 12000
rect 14348 11940 14352 11996
rect 14352 11940 14408 11996
rect 14408 11940 14412 11996
rect 14348 11936 14412 11940
rect 14428 11996 14492 12000
rect 14428 11940 14432 11996
rect 14432 11940 14488 11996
rect 14488 11940 14492 11996
rect 14428 11936 14492 11940
rect 14508 11996 14572 12000
rect 14508 11940 14512 11996
rect 14512 11940 14568 11996
rect 14568 11940 14572 11996
rect 14508 11936 14572 11940
rect 18707 11996 18771 12000
rect 18707 11940 18711 11996
rect 18711 11940 18767 11996
rect 18767 11940 18771 11996
rect 18707 11936 18771 11940
rect 18787 11996 18851 12000
rect 18787 11940 18791 11996
rect 18791 11940 18847 11996
rect 18847 11940 18851 11996
rect 18787 11936 18851 11940
rect 18867 11996 18931 12000
rect 18867 11940 18871 11996
rect 18871 11940 18927 11996
rect 18927 11940 18931 11996
rect 18867 11936 18931 11940
rect 18947 11996 19011 12000
rect 18947 11940 18951 11996
rect 18951 11940 19007 11996
rect 19007 11940 19011 11996
rect 18947 11936 19011 11940
rect 13860 11928 13924 11932
rect 13860 11872 13874 11928
rect 13874 11872 13924 11928
rect 13860 11868 13924 11872
rect 3171 11452 3235 11456
rect 3171 11396 3175 11452
rect 3175 11396 3231 11452
rect 3231 11396 3235 11452
rect 3171 11392 3235 11396
rect 3251 11452 3315 11456
rect 3251 11396 3255 11452
rect 3255 11396 3311 11452
rect 3311 11396 3315 11452
rect 3251 11392 3315 11396
rect 3331 11452 3395 11456
rect 3331 11396 3335 11452
rect 3335 11396 3391 11452
rect 3391 11396 3395 11452
rect 3331 11392 3395 11396
rect 3411 11452 3475 11456
rect 3411 11396 3415 11452
rect 3415 11396 3471 11452
rect 3471 11396 3475 11452
rect 3411 11392 3475 11396
rect 7610 11452 7674 11456
rect 7610 11396 7614 11452
rect 7614 11396 7670 11452
rect 7670 11396 7674 11452
rect 7610 11392 7674 11396
rect 7690 11452 7754 11456
rect 7690 11396 7694 11452
rect 7694 11396 7750 11452
rect 7750 11396 7754 11452
rect 7690 11392 7754 11396
rect 7770 11452 7834 11456
rect 7770 11396 7774 11452
rect 7774 11396 7830 11452
rect 7830 11396 7834 11452
rect 7770 11392 7834 11396
rect 7850 11452 7914 11456
rect 7850 11396 7854 11452
rect 7854 11396 7910 11452
rect 7910 11396 7914 11452
rect 7850 11392 7914 11396
rect 12049 11452 12113 11456
rect 12049 11396 12053 11452
rect 12053 11396 12109 11452
rect 12109 11396 12113 11452
rect 12049 11392 12113 11396
rect 12129 11452 12193 11456
rect 12129 11396 12133 11452
rect 12133 11396 12189 11452
rect 12189 11396 12193 11452
rect 12129 11392 12193 11396
rect 12209 11452 12273 11456
rect 12209 11396 12213 11452
rect 12213 11396 12269 11452
rect 12269 11396 12273 11452
rect 12209 11392 12273 11396
rect 12289 11452 12353 11456
rect 12289 11396 12293 11452
rect 12293 11396 12349 11452
rect 12349 11396 12353 11452
rect 12289 11392 12353 11396
rect 16488 11452 16552 11456
rect 16488 11396 16492 11452
rect 16492 11396 16548 11452
rect 16548 11396 16552 11452
rect 16488 11392 16552 11396
rect 16568 11452 16632 11456
rect 16568 11396 16572 11452
rect 16572 11396 16628 11452
rect 16628 11396 16632 11452
rect 16568 11392 16632 11396
rect 16648 11452 16712 11456
rect 16648 11396 16652 11452
rect 16652 11396 16708 11452
rect 16708 11396 16712 11452
rect 16648 11392 16712 11396
rect 16728 11452 16792 11456
rect 16728 11396 16732 11452
rect 16732 11396 16788 11452
rect 16788 11396 16792 11452
rect 16728 11392 16792 11396
rect 15700 11324 15764 11388
rect 16988 11052 17052 11116
rect 5390 10908 5454 10912
rect 5390 10852 5394 10908
rect 5394 10852 5450 10908
rect 5450 10852 5454 10908
rect 5390 10848 5454 10852
rect 5470 10908 5534 10912
rect 5470 10852 5474 10908
rect 5474 10852 5530 10908
rect 5530 10852 5534 10908
rect 5470 10848 5534 10852
rect 5550 10908 5614 10912
rect 5550 10852 5554 10908
rect 5554 10852 5610 10908
rect 5610 10852 5614 10908
rect 5550 10848 5614 10852
rect 5630 10908 5694 10912
rect 5630 10852 5634 10908
rect 5634 10852 5690 10908
rect 5690 10852 5694 10908
rect 5630 10848 5694 10852
rect 9829 10908 9893 10912
rect 9829 10852 9833 10908
rect 9833 10852 9889 10908
rect 9889 10852 9893 10908
rect 9829 10848 9893 10852
rect 9909 10908 9973 10912
rect 9909 10852 9913 10908
rect 9913 10852 9969 10908
rect 9969 10852 9973 10908
rect 9909 10848 9973 10852
rect 9989 10908 10053 10912
rect 9989 10852 9993 10908
rect 9993 10852 10049 10908
rect 10049 10852 10053 10908
rect 9989 10848 10053 10852
rect 10069 10908 10133 10912
rect 10069 10852 10073 10908
rect 10073 10852 10129 10908
rect 10129 10852 10133 10908
rect 10069 10848 10133 10852
rect 14268 10908 14332 10912
rect 14268 10852 14272 10908
rect 14272 10852 14328 10908
rect 14328 10852 14332 10908
rect 14268 10848 14332 10852
rect 14348 10908 14412 10912
rect 14348 10852 14352 10908
rect 14352 10852 14408 10908
rect 14408 10852 14412 10908
rect 14348 10848 14412 10852
rect 14428 10908 14492 10912
rect 14428 10852 14432 10908
rect 14432 10852 14488 10908
rect 14488 10852 14492 10908
rect 14428 10848 14492 10852
rect 14508 10908 14572 10912
rect 14508 10852 14512 10908
rect 14512 10852 14568 10908
rect 14568 10852 14572 10908
rect 14508 10848 14572 10852
rect 18707 10908 18771 10912
rect 18707 10852 18711 10908
rect 18711 10852 18767 10908
rect 18767 10852 18771 10908
rect 18707 10848 18771 10852
rect 18787 10908 18851 10912
rect 18787 10852 18791 10908
rect 18791 10852 18847 10908
rect 18847 10852 18851 10908
rect 18787 10848 18851 10852
rect 18867 10908 18931 10912
rect 18867 10852 18871 10908
rect 18871 10852 18927 10908
rect 18927 10852 18931 10908
rect 18867 10848 18931 10852
rect 18947 10908 19011 10912
rect 18947 10852 18951 10908
rect 18951 10852 19007 10908
rect 19007 10852 19011 10908
rect 18947 10848 19011 10852
rect 3171 10364 3235 10368
rect 3171 10308 3175 10364
rect 3175 10308 3231 10364
rect 3231 10308 3235 10364
rect 3171 10304 3235 10308
rect 3251 10364 3315 10368
rect 3251 10308 3255 10364
rect 3255 10308 3311 10364
rect 3311 10308 3315 10364
rect 3251 10304 3315 10308
rect 3331 10364 3395 10368
rect 3331 10308 3335 10364
rect 3335 10308 3391 10364
rect 3391 10308 3395 10364
rect 3331 10304 3395 10308
rect 3411 10364 3475 10368
rect 3411 10308 3415 10364
rect 3415 10308 3471 10364
rect 3471 10308 3475 10364
rect 3411 10304 3475 10308
rect 7610 10364 7674 10368
rect 7610 10308 7614 10364
rect 7614 10308 7670 10364
rect 7670 10308 7674 10364
rect 7610 10304 7674 10308
rect 7690 10364 7754 10368
rect 7690 10308 7694 10364
rect 7694 10308 7750 10364
rect 7750 10308 7754 10364
rect 7690 10304 7754 10308
rect 7770 10364 7834 10368
rect 7770 10308 7774 10364
rect 7774 10308 7830 10364
rect 7830 10308 7834 10364
rect 7770 10304 7834 10308
rect 7850 10364 7914 10368
rect 7850 10308 7854 10364
rect 7854 10308 7910 10364
rect 7910 10308 7914 10364
rect 7850 10304 7914 10308
rect 12049 10364 12113 10368
rect 12049 10308 12053 10364
rect 12053 10308 12109 10364
rect 12109 10308 12113 10364
rect 12049 10304 12113 10308
rect 12129 10364 12193 10368
rect 12129 10308 12133 10364
rect 12133 10308 12189 10364
rect 12189 10308 12193 10364
rect 12129 10304 12193 10308
rect 12209 10364 12273 10368
rect 12209 10308 12213 10364
rect 12213 10308 12269 10364
rect 12269 10308 12273 10364
rect 12209 10304 12273 10308
rect 12289 10364 12353 10368
rect 12289 10308 12293 10364
rect 12293 10308 12349 10364
rect 12349 10308 12353 10364
rect 12289 10304 12353 10308
rect 16488 10364 16552 10368
rect 16488 10308 16492 10364
rect 16492 10308 16548 10364
rect 16548 10308 16552 10364
rect 16488 10304 16552 10308
rect 16568 10364 16632 10368
rect 16568 10308 16572 10364
rect 16572 10308 16628 10364
rect 16628 10308 16632 10364
rect 16568 10304 16632 10308
rect 16648 10364 16712 10368
rect 16648 10308 16652 10364
rect 16652 10308 16708 10364
rect 16708 10308 16712 10364
rect 16648 10304 16712 10308
rect 16728 10364 16792 10368
rect 16728 10308 16732 10364
rect 16732 10308 16788 10364
rect 16788 10308 16792 10364
rect 16728 10304 16792 10308
rect 5390 9820 5454 9824
rect 5390 9764 5394 9820
rect 5394 9764 5450 9820
rect 5450 9764 5454 9820
rect 5390 9760 5454 9764
rect 5470 9820 5534 9824
rect 5470 9764 5474 9820
rect 5474 9764 5530 9820
rect 5530 9764 5534 9820
rect 5470 9760 5534 9764
rect 5550 9820 5614 9824
rect 5550 9764 5554 9820
rect 5554 9764 5610 9820
rect 5610 9764 5614 9820
rect 5550 9760 5614 9764
rect 5630 9820 5694 9824
rect 5630 9764 5634 9820
rect 5634 9764 5690 9820
rect 5690 9764 5694 9820
rect 5630 9760 5694 9764
rect 9829 9820 9893 9824
rect 9829 9764 9833 9820
rect 9833 9764 9889 9820
rect 9889 9764 9893 9820
rect 9829 9760 9893 9764
rect 9909 9820 9973 9824
rect 9909 9764 9913 9820
rect 9913 9764 9969 9820
rect 9969 9764 9973 9820
rect 9909 9760 9973 9764
rect 9989 9820 10053 9824
rect 9989 9764 9993 9820
rect 9993 9764 10049 9820
rect 10049 9764 10053 9820
rect 9989 9760 10053 9764
rect 10069 9820 10133 9824
rect 10069 9764 10073 9820
rect 10073 9764 10129 9820
rect 10129 9764 10133 9820
rect 10069 9760 10133 9764
rect 14268 9820 14332 9824
rect 14268 9764 14272 9820
rect 14272 9764 14328 9820
rect 14328 9764 14332 9820
rect 14268 9760 14332 9764
rect 14348 9820 14412 9824
rect 14348 9764 14352 9820
rect 14352 9764 14408 9820
rect 14408 9764 14412 9820
rect 14348 9760 14412 9764
rect 14428 9820 14492 9824
rect 14428 9764 14432 9820
rect 14432 9764 14488 9820
rect 14488 9764 14492 9820
rect 14428 9760 14492 9764
rect 14508 9820 14572 9824
rect 14508 9764 14512 9820
rect 14512 9764 14568 9820
rect 14568 9764 14572 9820
rect 14508 9760 14572 9764
rect 18707 9820 18771 9824
rect 18707 9764 18711 9820
rect 18711 9764 18767 9820
rect 18767 9764 18771 9820
rect 18707 9760 18771 9764
rect 18787 9820 18851 9824
rect 18787 9764 18791 9820
rect 18791 9764 18847 9820
rect 18847 9764 18851 9820
rect 18787 9760 18851 9764
rect 18867 9820 18931 9824
rect 18867 9764 18871 9820
rect 18871 9764 18927 9820
rect 18927 9764 18931 9820
rect 18867 9760 18931 9764
rect 18947 9820 19011 9824
rect 18947 9764 18951 9820
rect 18951 9764 19007 9820
rect 19007 9764 19011 9820
rect 18947 9760 19011 9764
rect 3171 9276 3235 9280
rect 3171 9220 3175 9276
rect 3175 9220 3231 9276
rect 3231 9220 3235 9276
rect 3171 9216 3235 9220
rect 3251 9276 3315 9280
rect 3251 9220 3255 9276
rect 3255 9220 3311 9276
rect 3311 9220 3315 9276
rect 3251 9216 3315 9220
rect 3331 9276 3395 9280
rect 3331 9220 3335 9276
rect 3335 9220 3391 9276
rect 3391 9220 3395 9276
rect 3331 9216 3395 9220
rect 3411 9276 3475 9280
rect 3411 9220 3415 9276
rect 3415 9220 3471 9276
rect 3471 9220 3475 9276
rect 3411 9216 3475 9220
rect 7610 9276 7674 9280
rect 7610 9220 7614 9276
rect 7614 9220 7670 9276
rect 7670 9220 7674 9276
rect 7610 9216 7674 9220
rect 7690 9276 7754 9280
rect 7690 9220 7694 9276
rect 7694 9220 7750 9276
rect 7750 9220 7754 9276
rect 7690 9216 7754 9220
rect 7770 9276 7834 9280
rect 7770 9220 7774 9276
rect 7774 9220 7830 9276
rect 7830 9220 7834 9276
rect 7770 9216 7834 9220
rect 7850 9276 7914 9280
rect 7850 9220 7854 9276
rect 7854 9220 7910 9276
rect 7910 9220 7914 9276
rect 7850 9216 7914 9220
rect 12049 9276 12113 9280
rect 12049 9220 12053 9276
rect 12053 9220 12109 9276
rect 12109 9220 12113 9276
rect 12049 9216 12113 9220
rect 12129 9276 12193 9280
rect 12129 9220 12133 9276
rect 12133 9220 12189 9276
rect 12189 9220 12193 9276
rect 12129 9216 12193 9220
rect 12209 9276 12273 9280
rect 12209 9220 12213 9276
rect 12213 9220 12269 9276
rect 12269 9220 12273 9276
rect 12209 9216 12273 9220
rect 12289 9276 12353 9280
rect 12289 9220 12293 9276
rect 12293 9220 12349 9276
rect 12349 9220 12353 9276
rect 12289 9216 12353 9220
rect 16488 9276 16552 9280
rect 16488 9220 16492 9276
rect 16492 9220 16548 9276
rect 16548 9220 16552 9276
rect 16488 9216 16552 9220
rect 16568 9276 16632 9280
rect 16568 9220 16572 9276
rect 16572 9220 16628 9276
rect 16628 9220 16632 9276
rect 16568 9216 16632 9220
rect 16648 9276 16712 9280
rect 16648 9220 16652 9276
rect 16652 9220 16708 9276
rect 16708 9220 16712 9276
rect 16648 9216 16712 9220
rect 16728 9276 16792 9280
rect 16728 9220 16732 9276
rect 16732 9220 16788 9276
rect 16788 9220 16792 9276
rect 16728 9216 16792 9220
rect 5390 8732 5454 8736
rect 5390 8676 5394 8732
rect 5394 8676 5450 8732
rect 5450 8676 5454 8732
rect 5390 8672 5454 8676
rect 5470 8732 5534 8736
rect 5470 8676 5474 8732
rect 5474 8676 5530 8732
rect 5530 8676 5534 8732
rect 5470 8672 5534 8676
rect 5550 8732 5614 8736
rect 5550 8676 5554 8732
rect 5554 8676 5610 8732
rect 5610 8676 5614 8732
rect 5550 8672 5614 8676
rect 5630 8732 5694 8736
rect 5630 8676 5634 8732
rect 5634 8676 5690 8732
rect 5690 8676 5694 8732
rect 5630 8672 5694 8676
rect 9829 8732 9893 8736
rect 9829 8676 9833 8732
rect 9833 8676 9889 8732
rect 9889 8676 9893 8732
rect 9829 8672 9893 8676
rect 9909 8732 9973 8736
rect 9909 8676 9913 8732
rect 9913 8676 9969 8732
rect 9969 8676 9973 8732
rect 9909 8672 9973 8676
rect 9989 8732 10053 8736
rect 9989 8676 9993 8732
rect 9993 8676 10049 8732
rect 10049 8676 10053 8732
rect 9989 8672 10053 8676
rect 10069 8732 10133 8736
rect 10069 8676 10073 8732
rect 10073 8676 10129 8732
rect 10129 8676 10133 8732
rect 10069 8672 10133 8676
rect 14268 8732 14332 8736
rect 14268 8676 14272 8732
rect 14272 8676 14328 8732
rect 14328 8676 14332 8732
rect 14268 8672 14332 8676
rect 14348 8732 14412 8736
rect 14348 8676 14352 8732
rect 14352 8676 14408 8732
rect 14408 8676 14412 8732
rect 14348 8672 14412 8676
rect 14428 8732 14492 8736
rect 14428 8676 14432 8732
rect 14432 8676 14488 8732
rect 14488 8676 14492 8732
rect 14428 8672 14492 8676
rect 14508 8732 14572 8736
rect 14508 8676 14512 8732
rect 14512 8676 14568 8732
rect 14568 8676 14572 8732
rect 14508 8672 14572 8676
rect 18707 8732 18771 8736
rect 18707 8676 18711 8732
rect 18711 8676 18767 8732
rect 18767 8676 18771 8732
rect 18707 8672 18771 8676
rect 18787 8732 18851 8736
rect 18787 8676 18791 8732
rect 18791 8676 18847 8732
rect 18847 8676 18851 8732
rect 18787 8672 18851 8676
rect 18867 8732 18931 8736
rect 18867 8676 18871 8732
rect 18871 8676 18927 8732
rect 18927 8676 18931 8732
rect 18867 8672 18931 8676
rect 18947 8732 19011 8736
rect 18947 8676 18951 8732
rect 18951 8676 19007 8732
rect 19007 8676 19011 8732
rect 18947 8672 19011 8676
rect 16252 8468 16316 8532
rect 3171 8188 3235 8192
rect 3171 8132 3175 8188
rect 3175 8132 3231 8188
rect 3231 8132 3235 8188
rect 3171 8128 3235 8132
rect 3251 8188 3315 8192
rect 3251 8132 3255 8188
rect 3255 8132 3311 8188
rect 3311 8132 3315 8188
rect 3251 8128 3315 8132
rect 3331 8188 3395 8192
rect 3331 8132 3335 8188
rect 3335 8132 3391 8188
rect 3391 8132 3395 8188
rect 3331 8128 3395 8132
rect 3411 8188 3475 8192
rect 3411 8132 3415 8188
rect 3415 8132 3471 8188
rect 3471 8132 3475 8188
rect 3411 8128 3475 8132
rect 7610 8188 7674 8192
rect 7610 8132 7614 8188
rect 7614 8132 7670 8188
rect 7670 8132 7674 8188
rect 7610 8128 7674 8132
rect 7690 8188 7754 8192
rect 7690 8132 7694 8188
rect 7694 8132 7750 8188
rect 7750 8132 7754 8188
rect 7690 8128 7754 8132
rect 7770 8188 7834 8192
rect 7770 8132 7774 8188
rect 7774 8132 7830 8188
rect 7830 8132 7834 8188
rect 7770 8128 7834 8132
rect 7850 8188 7914 8192
rect 7850 8132 7854 8188
rect 7854 8132 7910 8188
rect 7910 8132 7914 8188
rect 7850 8128 7914 8132
rect 12049 8188 12113 8192
rect 12049 8132 12053 8188
rect 12053 8132 12109 8188
rect 12109 8132 12113 8188
rect 12049 8128 12113 8132
rect 12129 8188 12193 8192
rect 12129 8132 12133 8188
rect 12133 8132 12189 8188
rect 12189 8132 12193 8188
rect 12129 8128 12193 8132
rect 12209 8188 12273 8192
rect 12209 8132 12213 8188
rect 12213 8132 12269 8188
rect 12269 8132 12273 8188
rect 12209 8128 12273 8132
rect 12289 8188 12353 8192
rect 12289 8132 12293 8188
rect 12293 8132 12349 8188
rect 12349 8132 12353 8188
rect 12289 8128 12353 8132
rect 16488 8188 16552 8192
rect 16488 8132 16492 8188
rect 16492 8132 16548 8188
rect 16548 8132 16552 8188
rect 16488 8128 16552 8132
rect 16568 8188 16632 8192
rect 16568 8132 16572 8188
rect 16572 8132 16628 8188
rect 16628 8132 16632 8188
rect 16568 8128 16632 8132
rect 16648 8188 16712 8192
rect 16648 8132 16652 8188
rect 16652 8132 16708 8188
rect 16708 8132 16712 8188
rect 16648 8128 16712 8132
rect 16728 8188 16792 8192
rect 16728 8132 16732 8188
rect 16732 8132 16788 8188
rect 16788 8132 16792 8188
rect 16728 8128 16792 8132
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 16251 18596 16317 18597
rect 16251 18532 16252 18596
rect 16316 18532 16317 18596
rect 16251 18531 16317 18532
rect 3163 16896 3483 17456
rect 3163 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3483 16896
rect 3163 15808 3483 16832
rect 3163 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3483 15808
rect 3163 14720 3483 15744
rect 3163 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3483 14720
rect 3163 13632 3483 14656
rect 3163 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3483 13632
rect 3163 12544 3483 13568
rect 3163 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3483 12544
rect 3163 11456 3483 12480
rect 3163 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3483 11456
rect 3163 10368 3483 11392
rect 3163 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3483 10368
rect 3163 9280 3483 10304
rect 3163 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3483 9280
rect 3163 8192 3483 9216
rect 3163 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3483 8192
rect 3163 7104 3483 8128
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 17440 5702 17456
rect 5382 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5702 17440
rect 5382 16352 5702 17376
rect 5382 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5702 16352
rect 5382 15264 5702 16288
rect 5382 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5702 15264
rect 5382 14176 5702 15200
rect 5382 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5702 14176
rect 5382 13088 5702 14112
rect 5382 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5702 13088
rect 5382 12000 5702 13024
rect 5382 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5702 12000
rect 5382 10912 5702 11936
rect 5382 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5702 10912
rect 5382 9824 5702 10848
rect 5382 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5702 9824
rect 5382 8736 5702 9760
rect 5382 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5702 8736
rect 5382 7648 5702 8672
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 16896 7922 17456
rect 7602 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7922 16896
rect 7602 15808 7922 16832
rect 7602 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7922 15808
rect 7602 14720 7922 15744
rect 7602 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7922 14720
rect 7602 13632 7922 14656
rect 7602 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7922 13632
rect 7602 12544 7922 13568
rect 7602 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7922 12544
rect 7602 11456 7922 12480
rect 7602 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7922 11456
rect 7602 10368 7922 11392
rect 7602 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7922 10368
rect 7602 9280 7922 10304
rect 7602 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7922 9280
rect 7602 8192 7922 9216
rect 7602 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7922 8192
rect 7602 7104 7922 8128
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 17440 10141 17456
rect 9821 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10141 17440
rect 9821 16352 10141 17376
rect 9821 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10141 16352
rect 9821 15264 10141 16288
rect 12041 16896 12361 17456
rect 12041 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12361 16896
rect 10547 16148 10613 16149
rect 10547 16084 10548 16148
rect 10612 16084 10613 16148
rect 10547 16083 10613 16084
rect 9821 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10141 15264
rect 9821 14176 10141 15200
rect 9821 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10141 14176
rect 9821 13088 10141 14112
rect 9821 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10141 13088
rect 9821 12000 10141 13024
rect 10550 12885 10610 16083
rect 12041 15808 12361 16832
rect 12041 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12361 15808
rect 11099 15604 11165 15605
rect 11099 15540 11100 15604
rect 11164 15540 11165 15604
rect 11099 15539 11165 15540
rect 11102 14109 11162 15539
rect 12041 14720 12361 15744
rect 14260 17440 14580 17456
rect 14260 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14580 17440
rect 14260 16352 14580 17376
rect 14260 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14580 16352
rect 13859 15604 13925 15605
rect 13859 15540 13860 15604
rect 13924 15540 13925 15604
rect 13859 15539 13925 15540
rect 12041 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12361 14720
rect 11099 14108 11165 14109
rect 11099 14044 11100 14108
rect 11164 14044 11165 14108
rect 11099 14043 11165 14044
rect 12041 13632 12361 14656
rect 12939 14516 13005 14517
rect 12939 14452 12940 14516
rect 13004 14452 13005 14516
rect 12939 14451 13005 14452
rect 12942 13701 13002 14451
rect 12939 13700 13005 13701
rect 12939 13636 12940 13700
rect 13004 13636 13005 13700
rect 12939 13635 13005 13636
rect 12041 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12361 13632
rect 10547 12884 10613 12885
rect 10547 12820 10548 12884
rect 10612 12820 10613 12884
rect 10547 12819 10613 12820
rect 9821 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10141 12000
rect 9821 10912 10141 11936
rect 9821 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10141 10912
rect 9821 9824 10141 10848
rect 9821 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10141 9824
rect 9821 8736 10141 9760
rect 9821 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10141 8736
rect 9821 7648 10141 8672
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 12544 12361 13568
rect 12041 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12361 12544
rect 12041 11456 12361 12480
rect 13862 11933 13922 15539
rect 14260 15264 14580 16288
rect 15883 16284 15949 16285
rect 15883 16220 15884 16284
rect 15948 16220 15949 16284
rect 15883 16219 15949 16220
rect 14260 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14580 15264
rect 14260 14176 14580 15200
rect 14260 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14580 14176
rect 14260 13088 14580 14112
rect 15699 13836 15765 13837
rect 15699 13772 15700 13836
rect 15764 13772 15765 13836
rect 15699 13771 15765 13772
rect 14260 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14580 13088
rect 14260 12000 14580 13024
rect 14260 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14580 12000
rect 13859 11932 13925 11933
rect 13859 11868 13860 11932
rect 13924 11868 13925 11932
rect 13859 11867 13925 11868
rect 12041 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12361 11456
rect 12041 10368 12361 11392
rect 12041 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12361 10368
rect 12041 9280 12361 10304
rect 12041 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12361 9280
rect 12041 8192 12361 9216
rect 12041 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12361 8192
rect 12041 7104 12361 8128
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 10912 14580 11936
rect 15702 11389 15762 13771
rect 15886 12069 15946 16219
rect 16067 14516 16133 14517
rect 16067 14452 16068 14516
rect 16132 14452 16133 14516
rect 16067 14451 16133 14452
rect 16070 12477 16130 14451
rect 16067 12476 16133 12477
rect 16067 12412 16068 12476
rect 16132 12412 16133 12476
rect 16067 12411 16133 12412
rect 15883 12068 15949 12069
rect 15883 12004 15884 12068
rect 15948 12004 15949 12068
rect 15883 12003 15949 12004
rect 15699 11388 15765 11389
rect 15699 11324 15700 11388
rect 15764 11324 15765 11388
rect 15699 11323 15765 11324
rect 14260 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14580 10912
rect 14260 9824 14580 10848
rect 14260 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14580 9824
rect 14260 8736 14580 9760
rect 14260 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14580 8736
rect 14260 7648 14580 8672
rect 16254 8533 16314 18531
rect 16480 16896 16800 17456
rect 16480 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16800 16896
rect 16480 15808 16800 16832
rect 16480 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16800 15808
rect 16480 14720 16800 15744
rect 16480 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16800 14720
rect 16480 13632 16800 14656
rect 16480 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16800 13632
rect 16480 12544 16800 13568
rect 18699 17440 19019 17456
rect 18699 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19019 17440
rect 18699 16352 19019 17376
rect 18699 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19019 16352
rect 18699 15264 19019 16288
rect 18699 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19019 15264
rect 18699 14176 19019 15200
rect 18699 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19019 14176
rect 16987 13292 17053 13293
rect 16987 13228 16988 13292
rect 17052 13228 17053 13292
rect 16987 13227 17053 13228
rect 16480 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16800 12544
rect 16480 11456 16800 12480
rect 16480 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16800 11456
rect 16480 10368 16800 11392
rect 16990 11117 17050 13227
rect 18699 13088 19019 14112
rect 18699 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19019 13088
rect 18699 12000 19019 13024
rect 18699 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19019 12000
rect 16987 11116 17053 11117
rect 16987 11052 16988 11116
rect 17052 11052 17053 11116
rect 16987 11051 17053 11052
rect 16480 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16800 10368
rect 16480 9280 16800 10304
rect 16480 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16800 9280
rect 16251 8532 16317 8533
rect 16251 8468 16252 8532
rect 16316 8468 16317 8532
rect 16251 8467 16317 8468
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 8192 16800 9216
rect 16480 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16800 8192
rect 16480 7104 16800 8128
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 10912 19019 11936
rect 18699 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19019 10912
rect 18699 9824 19019 10848
rect 18699 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19019 9824
rect 18699 8736 19019 9760
rect 18699 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19019 8736
rect 18699 7648 19019 8672
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout13_A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6808 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 17756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1666464484
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1666464484
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1666464484
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1666464484
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1666464484
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1666464484
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1666464484
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1666464484
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1666464484
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1666464484
transform 1 0 18400 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_8
timestamp 1666464484
transform 1 0 1840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1666464484
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1666464484
transform 1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1666464484
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_32
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1666464484
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_8
timestamp 1666464484
transform 1 0 1840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1666464484
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_188
timestamp 1666464484
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1666464484
transform 1 0 18400 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_8
timestamp 1666464484
transform 1 0 1840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1666464484
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1666464484
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_8
timestamp 1666464484
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1666464484
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1666464484
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1666464484
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1666464484
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1666464484
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1666464484
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1666464484
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1666464484
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_8
timestamp 1666464484
transform 1 0 1840 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_20
timestamp 1666464484
transform 1 0 2944 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_32
timestamp 1666464484
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1666464484
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1666464484
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1666464484
transform 1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_8
timestamp 1666464484
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1666464484
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_161
timestamp 1666464484
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1666464484
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1666464484
transform 1 0 17112 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_181
timestamp 1666464484
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1666464484
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1666464484
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1666464484
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_159
timestamp 1666464484
transform 1 0 15732 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1666464484
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1666464484
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1666464484
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1666464484
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1666464484
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1666464484
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_164
timestamp 1666464484
transform 1 0 16192 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_170
timestamp 1666464484
transform 1 0 16744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1666464484
transform 1 0 17112 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1666464484
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1666464484
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_8
timestamp 1666464484
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_20
timestamp 1666464484
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_32
timestamp 1666464484
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1666464484
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 1666464484
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1666464484
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1666464484
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1666464484
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1666464484
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1666464484
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1666464484
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1666464484
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_168
timestamp 1666464484
transform 1 0 16560 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_176
timestamp 1666464484
transform 1 0 17296 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_184
timestamp 1666464484
transform 1 0 18032 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1666464484
transform 1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1666464484
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1666464484
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1666464484
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_121
timestamp 1666464484
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1666464484
transform 1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1666464484
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1666464484
transform 1 0 14536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_157
timestamp 1666464484
transform 1 0 15548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1666464484
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1666464484
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1666464484
transform 1 0 18400 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_8
timestamp 1666464484
transform 1 0 1840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1666464484
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1666464484
transform 1 0 11960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1666464484
transform 1 0 12788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1666464484
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1666464484
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_166
timestamp 1666464484
transform 1 0 16376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1666464484
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_184
timestamp 1666464484
transform 1 0 18032 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_8
timestamp 1666464484
transform 1 0 1840 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_20
timestamp 1666464484
transform 1 0 2944 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_32
timestamp 1666464484
transform 1 0 4048 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_44
timestamp 1666464484
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_99
timestamp 1666464484
transform 1 0 10212 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1666464484
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1666464484
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1666464484
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_133
timestamp 1666464484
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_157
timestamp 1666464484
transform 1 0 15548 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1666464484
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_187
timestamp 1666464484
transform 1 0 18308 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1666464484
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1666464484
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1666464484
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_105
timestamp 1666464484
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1666464484
transform 1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1666464484
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1666464484
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1666464484
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1666464484
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1666464484
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_8
timestamp 1666464484
transform 1 0 1840 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_20
timestamp 1666464484
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_32
timestamp 1666464484
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1666464484
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_84
timestamp 1666464484
transform 1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_91
timestamp 1666464484
transform 1 0 9476 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_100
timestamp 1666464484
transform 1 0 10304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1666464484
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_129
timestamp 1666464484
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1666464484
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1666464484
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1666464484
transform 1 0 17572 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1666464484
transform 1 0 18400 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1666464484
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1666464484
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1666464484
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_75
timestamp 1666464484
transform 1 0 8004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1666464484
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1666464484
transform 1 0 9660 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1666464484
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_114
timestamp 1666464484
transform 1 0 11592 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1666464484
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1666464484
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1666464484
transform 1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_8
timestamp 1666464484
transform 1 0 1840 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_20
timestamp 1666464484
transform 1 0 2944 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_32
timestamp 1666464484
transform 1 0 4048 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_44
timestamp 1666464484
transform 1 0 5152 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1666464484
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 1666464484
transform 1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_87
timestamp 1666464484
transform 1 0 9108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_98
timestamp 1666464484
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1666464484
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1666464484
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1666464484
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1666464484
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_8
timestamp 1666464484
transform 1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 1666464484
transform 1 0 6256 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_63
timestamp 1666464484
transform 1 0 6900 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_72
timestamp 1666464484
transform 1 0 7728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1666464484
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_90
timestamp 1666464484
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1666464484
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1666464484
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_164
timestamp 1666464484
transform 1 0 16192 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp 1666464484
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_8
timestamp 1666464484
transform 1 0 1840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_22
timestamp 1666464484
transform 1 0 3128 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_34
timestamp 1666464484
transform 1 0 4232 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1666464484
transform 1 0 4968 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_47
timestamp 1666464484
transform 1 0 5428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1666464484
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_65
timestamp 1666464484
transform 1 0 7084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_75
timestamp 1666464484
transform 1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1666464484
transform 1 0 9016 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1666464484
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1666464484
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1666464484
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1666464484
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_8
timestamp 1666464484
transform 1 0 1840 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_16
timestamp 1666464484
transform 1 0 2576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_20
timestamp 1666464484
transform 1 0 2944 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_40
timestamp 1666464484
transform 1 0 4784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1666464484
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1666464484
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_63
timestamp 1666464484
transform 1 0 6900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_71
timestamp 1666464484
transform 1 0 7636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1666464484
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1666464484
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1666464484
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1666464484
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1666464484
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1666464484
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_187
timestamp 1666464484
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_8
timestamp 1666464484
transform 1 0 1840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_19
timestamp 1666464484
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1666464484
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_29
timestamp 1666464484
transform 1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_38
timestamp 1666464484
transform 1 0 4600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_46
timestamp 1666464484
transform 1 0 5336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1666464484
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_65
timestamp 1666464484
transform 1 0 7084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_73
timestamp 1666464484
transform 1 0 7820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_82
timestamp 1666464484
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1666464484
transform 1 0 8924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_89
timestamp 1666464484
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1666464484
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1666464484
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1666464484
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1666464484
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1666464484
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1666464484
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_188
timestamp 1666464484
transform 1 0 18400 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__or3b_1  _067_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _068_
timestamp 1666464484
transform -1 0 18216 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _069_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16560 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_2  _070_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _071_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17756 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _072_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _073_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _074_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17572 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _075_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14628 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _076_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16008 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _077_
timestamp 1666464484
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _078_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8648 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _079_
timestamp 1666464484
transform -1 0 17204 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _080_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7268 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _081_
timestamp 1666464484
transform -1 0 15180 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _082_
timestamp 1666464484
transform -1 0 17756 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _083_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9844 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _084_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _085_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9200 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _086_
timestamp 1666464484
transform -1 0 8648 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _087_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _088_
timestamp 1666464484
transform 1 0 14720 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _089_
timestamp 1666464484
transform 1 0 17848 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _090_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16376 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _091_
timestamp 1666464484
transform -1 0 5428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _092_
timestamp 1666464484
transform -1 0 15548 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _093_
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _094_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13800 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _095_
timestamp 1666464484
transform -1 0 17296 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _096_
timestamp 1666464484
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _097_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11684 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _098_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11960 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _099_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _100_
timestamp 1666464484
transform -1 0 10028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _101_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _102_
timestamp 1666464484
transform -1 0 18400 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _103_
timestamp 1666464484
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _104_
timestamp 1666464484
transform -1 0 16100 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _106_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _107_
timestamp 1666464484
transform -1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _108_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _109_
timestamp 1666464484
transform 1 0 8096 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _110_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1666464484
transform -1 0 14352 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _112_
timestamp 1666464484
transform 1 0 13156 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _113_
timestamp 1666464484
transform -1 0 6072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _114_
timestamp 1666464484
transform -1 0 12788 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _115_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11592 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _116_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12696 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _117_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8648 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _118_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8372 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _119_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _120_
timestamp 1666464484
transform -1 0 7084 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _121_
timestamp 1666464484
transform 1 0 9200 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _122_
timestamp 1666464484
transform -1 0 13524 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _123_
timestamp 1666464484
transform 1 0 6624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _124_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8004 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _125_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10672 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _126_
timestamp 1666464484
transform -1 0 10580 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _127_
timestamp 1666464484
transform -1 0 14536 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _128_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9384 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _129_
timestamp 1666464484
transform -1 0 11224 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _130_
timestamp 1666464484
transform 1 0 12696 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _131_
timestamp 1666464484
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _132_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12972 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1666464484
transform 1 0 18124 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _134_
timestamp 1666464484
transform 1 0 10948 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _135_
timestamp 1666464484
transform -1 0 12604 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1666464484
transform 1 0 18124 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _137_
timestamp 1666464484
transform -1 0 16376 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _138_
timestamp 1666464484
transform 1 0 9568 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _139_
timestamp 1666464484
transform 1 0 9476 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _140_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16468 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _141_
timestamp 1666464484
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _142_
timestamp 1666464484
transform 1 0 13340 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _143_
timestamp 1666464484
transform 1 0 11960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _144_
timestamp 1666464484
transform -1 0 13800 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _145_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16192 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _146_
timestamp 1666464484
transform 1 0 16560 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _147_
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _148_
timestamp 1666464484
transform 1 0 9384 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _149_
timestamp 1666464484
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _150_
timestamp 1666464484
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _151_
timestamp 1666464484
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _152_
timestamp 1666464484
transform 1 0 9752 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _153_
timestamp 1666464484
transform -1 0 16100 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _154_
timestamp 1666464484
transform -1 0 13800 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _155_
timestamp 1666464484
transform -1 0 14812 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _156_
timestamp 1666464484
transform -1 0 13800 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _157_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13340 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  fanout10 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15732 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout11 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1666464484
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1666464484
transform -1 0 7084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform 1 0 17480 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform 1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform 1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1666464484
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform -1 0 6072 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform 1 0 7268 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform -1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform -1 0 5336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_14 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_15
timestamp 1666464484
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_16
timestamp 1666464484
transform 1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_17
timestamp 1666464484
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_18
timestamp 1666464484
transform 1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_19
timestamp 1666464484
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_20
timestamp 1666464484
transform 1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_21
timestamp 1666464484
transform 1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_22
timestamp 1666464484
transform 1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_23
timestamp 1666464484
transform 1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_24
timestamp 1666464484
transform 1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_25
timestamp 1666464484
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_26
timestamp 1666464484
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_27
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_28
timestamp 1666464484
transform 1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_29
timestamp 1666464484
transform 1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_30
timestamp 1666464484
transform -1 0 16192 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_31
timestamp 1666464484
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_32
timestamp 1666464484
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_33
timestamp 1666464484
transform 1 0 4324 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_34
timestamp 1666464484
transform -1 0 7360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_35
timestamp 1666464484
transform 1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_36
timestamp 1666464484
transform -1 0 2944 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_37
timestamp 1666464484
transform -1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_38
timestamp 1666464484
transform -1 0 3128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_39
timestamp 1666464484
transform -1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_40
timestamp 1666464484
transform -1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_41
timestamp 1666464484
transform -1 0 1840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_42
timestamp 1666464484
transform -1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_43
timestamp 1666464484
transform -1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_44
timestamp 1666464484
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_45
timestamp 1666464484
transform -1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_46
timestamp 1666464484
transform -1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_47
timestamp 1666464484
transform -1 0 1840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_48
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_49
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_50
timestamp 1666464484
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_51
timestamp 1666464484
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_52
timestamp 1666464484
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_53
timestamp 1666464484
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_54
timestamp 1666464484
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_55
timestamp 1666464484
transform 1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_56
timestamp 1666464484
transform 1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_57
timestamp 1666464484
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_58
timestamp 1666464484
transform 1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_59
timestamp 1666464484
transform 1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_60
timestamp 1666464484
transform 1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_61
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_62
timestamp 1666464484
transform 1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_63
timestamp 1666464484
transform 1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_64
timestamp 1666464484
transform 1 0 12420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_65
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_66
timestamp 1666464484
transform 1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_67
timestamp 1666464484
transform 1 0 16192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_68
timestamp 1666464484
transform 1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_69
timestamp 1666464484
transform -1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_70
timestamp 1666464484
transform -1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_71
timestamp 1666464484
transform -1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_72
timestamp 1666464484
transform -1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_73
timestamp 1666464484
transform -1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_74
timestamp 1666464484
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_75
timestamp 1666464484
transform -1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_76
timestamp 1666464484
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_77
timestamp 1666464484
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_78
timestamp 1666464484
transform -1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_79
timestamp 1666464484
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_80
timestamp 1666464484
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_81
timestamp 1666464484
transform -1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_82
timestamp 1666464484
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_83
timestamp 1666464484
transform -1 0 2484 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal3 s 19200 960 20000 1080 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 19200 13200 20000 13320 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 19200 14424 20000 14544 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 19200 15648 20000 15768 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 19200 16872 20000 16992 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 19200 18096 20000 18216 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 19522 19200 19578 20000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 17314 19200 17370 20000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 15106 19200 15162 20000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 12898 19200 12954 20000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 10690 19200 10746 20000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 19200 2184 20000 2304 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 8482 19200 8538 20000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 6274 19200 6330 20000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 4066 19200 4122 20000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 1858 19200 1914 20000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 19200 3408 20000 3528 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 19200 5856 20000 5976 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 19200 7080 20000 7200 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 19200 8304 20000 8424 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 19200 10752 20000 10872 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 19200 1776 20000 1896 0 FreeSans 480 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 19200 14016 20000 14136 0 FreeSans 480 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 19200 15240 20000 15360 0 FreeSans 480 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 19200 16464 20000 16584 0 FreeSans 480 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 19200 17688 20000 17808 0 FreeSans 480 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 19200 18912 20000 19032 0 FreeSans 480 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 18050 19200 18106 20000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 15842 19200 15898 20000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 13634 19200 13690 20000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 11426 19200 11482 20000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 9218 19200 9274 20000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 7010 19200 7066 20000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 4802 19200 4858 20000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 2594 19200 2650 20000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 386 19200 442 20000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 19200 4224 20000 4344 0 FreeSans 480 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 19200 6672 20000 6792 0 FreeSans 480 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 19200 7896 20000 8016 0 FreeSans 480 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 19200 9120 20000 9240 0 FreeSans 480 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 19200 11568 20000 11688 0 FreeSans 480 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 19200 12792 20000 12912 0 FreeSans 480 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 19200 14832 20000 14952 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 19200 17280 20000 17400 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 19200 18504 20000 18624 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 18786 19200 18842 20000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 16578 19200 16634 20000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 14370 19200 14426 20000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 12162 19200 12218 20000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 9954 19200 10010 20000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 19200 2592 20000 2712 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 7746 19200 7802 20000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 5538 19200 5594 20000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 3330 19200 3386 20000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 1122 19200 1178 20000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 19200 5040 20000 5160 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 19200 7488 20000 7608 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 19200 9936 20000 10056 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 19200 12384 20000 12504 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 3163 2128 3483 17456 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 7602 2128 7922 17456 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 12041 2128 12361 17456 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 16480 2128 16800 17456 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 5382 2128 5702 17456 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 9821 2128 10141 17456 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 14260 2128 14580 17456 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 18699 2128 19019 17456 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 9982 16864 9982 16864 0 vccd1
rlabel via1 10061 17408 10061 17408 0 vssd1
rlabel metal2 8602 15402 8602 15402 0 _000_
rlabel metal1 9890 15538 9890 15538 0 _001_
rlabel metal2 13294 12852 13294 12852 0 _002_
rlabel metal1 14030 15538 14030 15538 0 _003_
rlabel metal1 14720 15062 14720 15062 0 _004_
rlabel metal2 13478 16932 13478 16932 0 _005_
rlabel metal2 16790 16303 16790 16303 0 _006_
rlabel metal2 10534 15113 10534 15113 0 _007_
rlabel metal2 7498 14824 7498 14824 0 _008_
rlabel metal1 10994 14518 10994 14518 0 _009_
rlabel metal1 13708 14314 13708 14314 0 _010_
rlabel metal1 15778 12274 15778 12274 0 _011_
rlabel metal1 13156 13362 13156 13362 0 _012_
rlabel metal1 12972 12886 12972 12886 0 _013_
rlabel metal2 15594 14790 15594 14790 0 _014_
rlabel metal1 14628 14450 14628 14450 0 _015_
rlabel metal2 11638 14467 11638 14467 0 _016_
rlabel metal1 13616 12342 13616 12342 0 _017_
rlabel metal2 6670 15844 6670 15844 0 _018_
rlabel metal1 10626 13702 10626 13702 0 _019_
rlabel metal2 12834 14926 12834 14926 0 _020_
rlabel metal1 12466 15980 12466 15980 0 _021_
rlabel metal1 13202 15946 13202 15946 0 _022_
rlabel metal2 11546 14722 11546 14722 0 _023_
rlabel metal2 12558 15504 12558 15504 0 _024_
rlabel metal1 16100 12682 16100 12682 0 _025_
rlabel metal1 9706 14926 9706 14926 0 _026_
rlabel metal2 17434 13702 17434 13702 0 _027_
rlabel metal1 17572 13498 17572 13498 0 _028_
rlabel metal1 16514 14926 16514 14926 0 _029_
rlabel metal2 16882 16745 16882 16745 0 _030_
rlabel metal1 16008 14042 16008 14042 0 _031_
rlabel metal1 8602 16490 8602 16490 0 _032_
rlabel metal1 16238 10778 16238 10778 0 _033_
rlabel metal1 7222 15470 7222 15470 0 _034_
rlabel metal2 16514 13209 16514 13209 0 _035_
rlabel metal1 16054 12240 16054 12240 0 _036_
rlabel metal1 10304 13702 10304 13702 0 _037_
rlabel metal2 15870 13855 15870 13855 0 _038_
rlabel metal1 8970 14246 8970 14246 0 _039_
rlabel metal2 16146 11951 16146 11951 0 _040_
rlabel metal1 17480 10778 17480 10778 0 _041_
rlabel metal2 15134 11526 15134 11526 0 _042_
rlabel metal2 16284 12716 16284 12716 0 _043_
rlabel via2 13386 13379 13386 13379 0 _044_
rlabel metal1 13616 11526 13616 11526 0 _045_
rlabel metal1 13432 13294 13432 13294 0 _046_
rlabel metal1 15778 13872 15778 13872 0 _047_
rlabel metal2 11178 14042 11178 14042 0 _048_
rlabel metal2 11822 12954 11822 12954 0 _049_
rlabel metal1 10902 13430 10902 13430 0 _050_
rlabel metal2 16238 14076 16238 14076 0 _051_
rlabel metal2 17940 12716 17940 12716 0 _052_
rlabel metal1 12788 11322 12788 11322 0 _053_
rlabel metal1 12282 12818 12282 12818 0 _054_
rlabel metal2 12742 14195 12742 14195 0 _055_
rlabel metal1 13754 11730 13754 11730 0 _056_
rlabel metal1 13018 14042 13018 14042 0 _057_
rlabel metal2 8878 15164 8878 15164 0 _058_
rlabel metal2 14214 11492 14214 11492 0 _059_
rlabel metal2 6026 14382 6026 14382 0 _060_
rlabel metal1 11868 12410 11868 12410 0 _061_
rlabel metal2 11914 14110 11914 14110 0 _062_
rlabel metal2 8418 13770 8418 13770 0 _063_
rlabel metal2 18078 14365 18078 14365 0 _064_
rlabel metal1 6670 15504 6670 15504 0 _065_
rlabel metal2 8234 15198 8234 15198 0 _066_
rlabel metal3 18362 13260 18362 13260 0 io_in[10]
rlabel metal1 18492 9554 18492 9554 0 io_in[8]
rlabel via2 18354 11747 18354 11747 0 io_in[9]
rlabel metal2 16836 19244 16836 19244 0 io_out[16]
rlabel metal2 14214 17663 14214 17663 0 io_out[17]
rlabel metal1 9752 17306 9752 17306 0 io_out[18]
rlabel metal2 9798 16779 9798 16779 0 io_out[19]
rlabel metal2 7958 16099 7958 16099 0 io_out[20]
rlabel metal1 5428 17306 5428 17306 0 io_out[21]
rlabel metal1 12029 12274 12029 12274 0 mod.cnter_enb_ovf_i1.cnt_val\[0\]
rlabel metal1 12742 12818 12742 12818 0 mod.cnter_enb_ovf_i1.cnt_val\[1\]
rlabel metal2 12650 12988 12650 12988 0 mod.cnter_enb_ovf_i1.cnt_val\[2\]
rlabel metal2 16330 13124 16330 13124 0 mod.cnter_enb_ovf_i1.cnt_val\[3\]
rlabel metal1 10074 14994 10074 14994 0 mod.cnter_enb_ovf_i1.cnt_val\[4\]
rlabel metal2 8694 15810 8694 15810 0 mod.cnter_enb_ovf_i1.overflow
rlabel metal1 8832 16082 8832 16082 0 mod.cnter_enb_ovf_i2.cnt_val\[0\]
rlabel metal2 7314 15045 7314 15045 0 mod.cnter_enb_ovf_i2.cnt_val\[1\]
rlabel metal2 6762 14382 6762 14382 0 mod.cnter_enb_ovf_i2.cnt_val\[2\]
rlabel metal1 13800 16422 13800 16422 0 mod.cnter_enb_ovf_i2.cnt_val\[3\]
rlabel metal1 8234 14314 8234 14314 0 mod.cnter_enb_ovf_i2.cnt_val\[4\]
rlabel metal1 14950 12206 14950 12206 0 mod.traffic_sm_inst.traffic_state\[0\]
rlabel metal1 17434 13736 17434 13736 0 mod.traffic_sm_inst.traffic_state\[1\]
rlabel metal1 15456 12206 15456 12206 0 mod.traffic_sm_inst.traffic_state\[2\]
rlabel metal1 14582 12410 14582 12410 0 mod.traffic_sm_inst.traffic_state\[3\]
rlabel metal2 17618 16592 17618 16592 0 mod.traffic_sm_inst.traffic_state\[4\]
rlabel metal1 17020 15946 17020 15946 0 mod.traffic_sm_inst.traffic_state\[5\]
rlabel metal1 16700 12818 16700 12818 0 mod.traffic_sm_inst.traffic_state\[6\]
rlabel metal2 17526 10438 17526 10438 0 net1
rlabel metal2 17342 15946 17342 15946 0 net10
rlabel metal2 17802 13600 17802 13600 0 net11
rlabel metal2 13754 17442 13754 17442 0 net12
rlabel metal2 6670 16728 6670 16728 0 net13
rlabel metal2 18354 2125 18354 2125 0 net14
rlabel metal2 18354 3281 18354 3281 0 net15
rlabel metal1 18768 4590 18768 4590 0 net16
rlabel via2 18354 5661 18354 5661 0 net17
rlabel via2 18354 6749 18354 6749 0 net18
rlabel via2 18354 7939 18354 7939 0 net19
rlabel metal1 12512 9418 12512 9418 0 net2
rlabel metal2 18354 8823 18354 8823 0 net20
rlabel metal2 17066 10319 17066 10319 0 net21
rlabel metal2 18354 11475 18354 11475 0 net22
rlabel via2 17733 12580 17733 12580 0 net23
rlabel metal1 18078 9486 18078 9486 0 net24
rlabel metal1 16330 9588 16330 9588 0 net25
rlabel metal3 17020 16320 17020 16320 0 net26
rlabel metal2 16054 16388 16054 16388 0 net27
rlabel metal2 15686 16932 15686 16932 0 net28
rlabel metal2 18124 15844 18124 15844 0 net29
rlabel metal2 18170 12036 18170 12036 0 net3
rlabel metal2 15916 17884 15916 17884 0 net30
rlabel metal2 13662 18370 13662 18370 0 net31
rlabel metal1 10304 15674 10304 15674 0 net32
rlabel metal1 6900 17034 6900 17034 0 net33
rlabel metal1 7084 14586 7084 14586 0 net34
rlabel metal1 4140 17170 4140 17170 0 net35
rlabel metal1 2668 16762 2668 16762 0 net36
rlabel metal1 1334 16014 1334 16014 0 net37
rlabel metal2 2898 16779 2898 16779 0 net38
rlabel metal3 1142 16252 1142 16252 0 net39
rlabel metal1 15778 10166 15778 10166 0 net4
rlabel metal3 1142 15028 1142 15028 0 net40
rlabel metal3 1142 13804 1142 13804 0 net41
rlabel metal3 1142 12580 1142 12580 0 net42
rlabel metal3 1142 11356 1142 11356 0 net43
rlabel metal3 1142 10132 1142 10132 0 net44
rlabel metal3 1142 8908 1142 8908 0 net45
rlabel metal3 1142 7684 1142 7684 0 net46
rlabel metal3 1142 6460 1142 6460 0 net47
rlabel via2 1610 5219 1610 5219 0 net48
rlabel metal3 1142 4012 1142 4012 0 net49
rlabel metal1 7222 17102 7222 17102 0 net5
rlabel metal3 1142 2788 1142 2788 0 net50
rlabel metal3 1142 1564 1142 1564 0 net51
rlabel metal2 17710 1921 17710 1921 0 net52
rlabel metal3 18868 2652 18868 2652 0 net53
rlabel via2 18354 3893 18354 3893 0 net54
rlabel via2 18354 5083 18354 5083 0 net55
rlabel via2 18354 6307 18354 6307 0 net56
rlabel via2 18354 7395 18354 7395 0 net57
rlabel via2 17066 8925 17066 8925 0 net58
rlabel metal2 17710 9775 17710 9775 0 net59
rlabel metal1 7452 17170 7452 17170 0 net6
rlabel metal2 18354 10727 18354 10727 0 net60
rlabel metal3 18914 12444 18914 12444 0 net61
rlabel metal3 18960 13668 18960 13668 0 net62
rlabel metal3 18868 14892 18868 14892 0 net63
rlabel metal3 13018 12444 13018 12444 0 net64
rlabel metal2 6210 16728 6210 16728 0 net65
rlabel metal3 17833 18564 17833 18564 0 net66
rlabel metal2 19090 19244 19090 19244 0 net67
rlabel metal1 3082 17170 3082 17170 0 net68
rlabel metal1 1380 16082 1380 16082 0 net69
rlabel metal1 6578 16558 6578 16558 0 net7
rlabel metal2 2806 16779 2806 16779 0 net70
rlabel metal3 1050 16660 1050 16660 0 net71
rlabel metal1 1564 14994 1564 14994 0 net72
rlabel metal3 1142 14212 1142 14212 0 net73
rlabel metal3 1142 12988 1142 12988 0 net74
rlabel metal3 1142 11764 1142 11764 0 net75
rlabel metal3 1142 10540 1142 10540 0 net76
rlabel metal3 1142 9316 1142 9316 0 net77
rlabel metal3 1142 8092 1142 8092 0 net78
rlabel metal3 1142 6868 1142 6868 0 net79
rlabel metal2 17158 16388 17158 16388 0 net8
rlabel metal3 1142 5644 1142 5644 0 net80
rlabel metal3 1142 4420 1142 4420 0 net81
rlabel metal3 1142 3196 1142 3196 0 net82
rlabel metal3 1464 1972 1464 1972 0 net83
rlabel metal1 8464 15606 8464 15606 0 net9
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
