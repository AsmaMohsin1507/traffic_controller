// This is the unpowered netlist.
module tiny_user_project (io_in,
    io_oeb,
    io_out);
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire net15;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net16;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net17;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net53;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net54;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net55;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire \mod.cnter_enb_ovf_i1.cnt_val[0] ;
 wire \mod.cnter_enb_ovf_i1.cnt_val[1] ;
 wire \mod.cnter_enb_ovf_i1.cnt_val[2] ;
 wire \mod.cnter_enb_ovf_i1.cnt_val[3] ;
 wire \mod.cnter_enb_ovf_i1.cnt_val[4] ;
 wire \mod.cnter_enb_ovf_i1.overflow ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[0] ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[1] ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[2] ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[3] ;
 wire \mod.cnter_enb_ovf_i2.cnt_val[4] ;
 wire \mod.traffic_sm_inst.traffic_state[0] ;
 wire \mod.traffic_sm_inst.traffic_state[1] ;
 wire \mod.traffic_sm_inst.traffic_state[2] ;
 wire \mod.traffic_sm_inst.traffic_state[3] ;
 wire \mod.traffic_sm_inst.traffic_state[4] ;
 wire \mod.traffic_sm_inst.traffic_state[5] ;
 wire \mod.traffic_sm_inst.traffic_state[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;

 sky130_fd_sc_hd__or3b_1 _067_ (.A(\mod.traffic_sm_inst.traffic_state[5] ),
    .B(\mod.traffic_sm_inst.traffic_state[4] ),
    .C_N(\mod.traffic_sm_inst.traffic_state[6] ),
    .X(_027_));
 sky130_fd_sc_hd__or3b_1 _068_ (.A(\mod.traffic_sm_inst.traffic_state[5] ),
    .B(\mod.traffic_sm_inst.traffic_state[6] ),
    .C_N(\mod.traffic_sm_inst.traffic_state[4] ),
    .X(_028_));
 sky130_fd_sc_hd__nor4_1 _069_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(\mod.traffic_sm_inst.traffic_state[1] ),
    .C(\mod.traffic_sm_inst.traffic_state[3] ),
    .D(\mod.traffic_sm_inst.traffic_state[2] ),
    .Y(_029_));
 sky130_fd_sc_hd__a21boi_2 _070_ (.A1(_027_),
    .A2(_028_),
    .B1_N(_029_),
    .Y(net8));
 sky130_fd_sc_hd__and4bb_1 _071_ (.A_N(\mod.traffic_sm_inst.traffic_state[4] ),
    .B_N(\mod.traffic_sm_inst.traffic_state[6] ),
    .C(_029_),
    .D(\mod.traffic_sm_inst.traffic_state[5] ),
    .X(_030_));
 sky130_fd_sc_hd__clkbuf_2 _072_ (.A(_030_),
    .X(net9));
 sky130_fd_sc_hd__nor2_1 _073_ (.A(net8),
    .B(net9),
    .Y(net7));
 sky130_fd_sc_hd__or4b_1 _074_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(\mod.traffic_sm_inst.traffic_state[1] ),
    .C(\mod.traffic_sm_inst.traffic_state[2] ),
    .D_N(\mod.traffic_sm_inst.traffic_state[3] ),
    .X(_031_));
 sky130_fd_sc_hd__or4b_2 _075_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(\mod.traffic_sm_inst.traffic_state[3] ),
    .C(\mod.traffic_sm_inst.traffic_state[2] ),
    .D_N(\mod.traffic_sm_inst.traffic_state[1] ),
    .X(_032_));
 sky130_fd_sc_hd__or3_1 _076_ (.A(\mod.traffic_sm_inst.traffic_state[5] ),
    .B(\mod.traffic_sm_inst.traffic_state[4] ),
    .C(\mod.traffic_sm_inst.traffic_state[6] ),
    .X(_033_));
 sky130_fd_sc_hd__clkbuf_2 _077_ (.A(_033_),
    .X(_034_));
 sky130_fd_sc_hd__a21oi_2 _078_ (.A1(_031_),
    .A2(_032_),
    .B1(_034_),
    .Y(net5));
 sky130_fd_sc_hd__or4b_1 _079_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(\mod.traffic_sm_inst.traffic_state[1] ),
    .C(\mod.traffic_sm_inst.traffic_state[3] ),
    .D_N(\mod.traffic_sm_inst.traffic_state[2] ),
    .X(_035_));
 sky130_fd_sc_hd__nor2_2 _080_ (.A(_034_),
    .B(_035_),
    .Y(net6));
 sky130_fd_sc_hd__nor2_1 _081_ (.A(net5),
    .B(net6),
    .Y(net4));
 sky130_fd_sc_hd__and4bb_1 _082_ (.A_N(\mod.traffic_sm_inst.traffic_state[5] ),
    .B_N(\mod.traffic_sm_inst.traffic_state[4] ),
    .C(\mod.traffic_sm_inst.traffic_state[6] ),
    .D(_029_),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _083_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .X(_037_));
 sky130_fd_sc_hd__and2b_1 _084_ (.A_N(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .X(_038_));
 sky130_fd_sc_hd__and3_1 _085_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .B(_037_),
    .C(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nor4_1 _086_ (.A(net8),
    .B(net9),
    .C(net5),
    .D(net6),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_1 _087_ (.A(\mod.traffic_sm_inst.traffic_state[0] ),
    .B(net1),
    .Y(_041_));
 sky130_fd_sc_hd__or3_1 _088_ (.A(\mod.traffic_sm_inst.traffic_state[1] ),
    .B(\mod.traffic_sm_inst.traffic_state[3] ),
    .C(\mod.traffic_sm_inst.traffic_state[2] ),
    .X(_042_));
 sky130_fd_sc_hd__or3_1 _089_ (.A(_034_),
    .B(_041_),
    .C(_042_),
    .X(_043_));
 sky130_fd_sc_hd__a22o_1 _090_ (.A1(_036_),
    .A2(_039_),
    .B1(_040_),
    .B2(_043_),
    .X(_011_));
 sky130_fd_sc_hd__nor2_1 _091_ (.A(_034_),
    .B(_032_),
    .Y(_044_));
 sky130_fd_sc_hd__or3b_1 _092_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .C_N(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .X(_045_));
 sky130_fd_sc_hd__or3_1 _093_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .C(_045_),
    .X(_046_));
 sky130_fd_sc_hd__a21bo_1 _094_ (.A1(_044_),
    .A2(_046_),
    .B1_N(_043_),
    .X(_012_));
 sky130_fd_sc_hd__and2b_1 _095_ (.A_N(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .B(_037_),
    .X(_047_));
 sky130_fd_sc_hd__a21bo_1 _096_ (.A1(_038_),
    .A2(_047_),
    .B1_N(net6),
    .X(_048_));
 sky130_fd_sc_hd__o31ai_1 _097_ (.A1(_034_),
    .A2(_032_),
    .A3(_046_),
    .B1(_048_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _098_ (.A(_045_),
    .Y(_049_));
 sky130_fd_sc_hd__nand3_1 _099_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .C(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__nor2_1 _100_ (.A(_034_),
    .B(_031_),
    .Y(_051_));
 sky130_fd_sc_hd__a32o_1 _101_ (.A1(net6),
    .A2(_038_),
    .A3(_047_),
    .B1(_050_),
    .B2(_051_),
    .X(_014_));
 sky130_fd_sc_hd__and3_1 _102_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .C(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .X(_052_));
 sky130_fd_sc_hd__nand2_1 _103_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .B(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__and4bb_1 _104_ (.A_N(\mod.traffic_sm_inst.traffic_state[5] ),
    .B_N(\mod.traffic_sm_inst.traffic_state[6] ),
    .C(_029_),
    .D(\mod.traffic_sm_inst.traffic_state[4] ),
    .X(_054_));
 sky130_fd_sc_hd__o21a_1 _105_ (.A1(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .A2(_053_),
    .B1(_054_),
    .X(_055_));
 sky130_fd_sc_hd__a41o_1 _106_ (.A1(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .A2(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .A3(_051_),
    .A4(_049_),
    .B1(_055_),
    .X(_015_));
 sky130_fd_sc_hd__nor2_1 _107_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .B(_053_),
    .Y(_056_));
 sky130_fd_sc_hd__and4b_1 _108_ (.A_N(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .C(_038_),
    .D(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .X(_057_));
 sky130_fd_sc_hd__and2b_1 _109_ (.A_N(_057_),
    .B(net9),
    .X(_058_));
 sky130_fd_sc_hd__a21o_1 _110_ (.A1(_054_),
    .A2(_056_),
    .B1(_058_),
    .X(_016_));
 sky130_fd_sc_hd__inv_2 _111_ (.A(_039_),
    .Y(_059_));
 sky130_fd_sc_hd__a22o_1 _112_ (.A1(_036_),
    .A2(_059_),
    .B1(_057_),
    .B2(net9),
    .X(_017_));
 sky130_fd_sc_hd__nor2_1 _113_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[3] ),
    .B(\mod.cnter_enb_ovf_i1.cnt_val[4] ),
    .Y(_060_));
 sky130_fd_sc_hd__and2_1 _114_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i1.cnt_val[0] ),
    .X(_061_));
 sky130_fd_sc_hd__o41a_1 _115_ (.A1(net8),
    .A2(net9),
    .A3(net5),
    .A4(net6),
    .B1(_061_),
    .X(_062_));
 sky130_fd_sc_hd__and3b_1 _116_ (.A_N(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .B(_060_),
    .C(_062_),
    .X(_063_));
 sky130_fd_sc_hd__clkbuf_1 _117_ (.A(_063_),
    .X(_000_));
 sky130_fd_sc_hd__xor2_1 _118_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .B(\mod.cnter_enb_ovf_i1.overflow ),
    .X(_006_));
 sky130_fd_sc_hd__a21oi_1 _119_ (.A1(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .A2(\mod.cnter_enb_ovf_i1.overflow ),
    .B1(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .Y(_064_));
 sky130_fd_sc_hd__and3_1 _120_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[1] ),
    .B(\mod.cnter_enb_ovf_i2.cnt_val[0] ),
    .C(\mod.cnter_enb_ovf_i1.overflow ),
    .X(_065_));
 sky130_fd_sc_hd__nor2_1 _121_ (.A(_064_),
    .B(_065_),
    .Y(_007_));
 sky130_fd_sc_hd__and2_1 _122_ (.A(\mod.cnter_enb_ovf_i1.overflow ),
    .B(_052_),
    .X(_066_));
 sky130_fd_sc_hd__nor2_1 _123_ (.A(\mod.cnter_enb_ovf_i2.cnt_val[2] ),
    .B(_065_),
    .Y(_018_));
 sky130_fd_sc_hd__a211oi_1 _124_ (.A1(\mod.cnter_enb_ovf_i1.overflow ),
    .A2(_039_),
    .B1(_066_),
    .C1(_018_),
    .Y(_008_));
 sky130_fd_sc_hd__a22oi_1 _125_ (.A1(\mod.cnter_enb_ovf_i1.overflow ),
    .A2(_039_),
    .B1(_066_),
    .B2(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .Y(_019_));
 sky130_fd_sc_hd__o21a_1 _126_ (.A1(\mod.cnter_enb_ovf_i2.cnt_val[3] ),
    .A2(_066_),
    .B1(_019_),
    .X(_009_));
 sky130_fd_sc_hd__a22o_1 _127_ (.A1(\mod.cnter_enb_ovf_i1.overflow ),
    .A2(_056_),
    .B1(_019_),
    .B2(\mod.cnter_enb_ovf_i2.cnt_val[4] ),
    .X(_010_));
 sky130_fd_sc_hd__xnor2_1 _128_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[0] ),
    .B(_040_),
    .Y(_001_));
 sky130_fd_sc_hd__o41a_1 _129_ (.A1(net8),
    .A2(net9),
    .A3(net5),
    .A4(net6),
    .B1(\mod.cnter_enb_ovf_i1.cnt_val[0] ),
    .X(_020_));
 sky130_fd_sc_hd__xor2_1 _130_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[1] ),
    .B(_020_),
    .X(_002_));
 sky130_fd_sc_hd__nor2_1 _131_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .B(_060_),
    .Y(_021_));
 sky130_fd_sc_hd__mux2_1 _132_ (.A0(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .A1(_021_),
    .S(_062_),
    .X(_022_));
 sky130_fd_sc_hd__clkbuf_1 _133_ (.A(_022_),
    .X(_003_));
 sky130_fd_sc_hd__xor2_1 _134_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[3] ),
    .B(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _135_ (.A0(\mod.cnter_enb_ovf_i1.cnt_val[3] ),
    .A1(_023_),
    .S(_062_),
    .X(_024_));
 sky130_fd_sc_hd__clkbuf_1 _136_ (.A(_024_),
    .X(_004_));
 sky130_fd_sc_hd__and3_1 _137_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[3] ),
    .B(\mod.cnter_enb_ovf_i1.cnt_val[2] ),
    .C(_061_),
    .X(_025_));
 sky130_fd_sc_hd__o41a_1 _138_ (.A1(net8),
    .A2(net9),
    .A3(net5),
    .A4(net6),
    .B1(_025_),
    .X(_026_));
 sky130_fd_sc_hd__xor2_1 _139_ (.A(\mod.cnter_enb_ovf_i1.cnt_val[4] ),
    .B(_026_),
    .X(_005_));
 sky130_fd_sc_hd__dfrtp_1 _140_ (.CLK(net12),
    .D(_006_),
    .RESET_B(net10),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[0] ));
 sky130_fd_sc_hd__dfrtp_1 _141_ (.CLK(net13),
    .D(_007_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[1] ));
 sky130_fd_sc_hd__dfrtp_1 _142_ (.CLK(net13),
    .D(_008_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[2] ));
 sky130_fd_sc_hd__dfrtp_1 _143_ (.CLK(net13),
    .D(_009_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[3] ));
 sky130_fd_sc_hd__dfrtp_1 _144_ (.CLK(net12),
    .D(_010_),
    .RESET_B(net10),
    .Q(\mod.cnter_enb_ovf_i2.cnt_val[4] ));
 sky130_fd_sc_hd__dfstp_1 _145_ (.CLK(net12),
    .D(_011_),
    .SET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _146_ (.CLK(net12),
    .D(_012_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _147_ (.CLK(net12),
    .D(_013_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _148_ (.CLK(net12),
    .D(_014_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _149_ (.CLK(net12),
    .D(_015_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _150_ (.CLK(net12),
    .D(_016_),
    .RESET_B(net10),
    .Q(\mod.traffic_sm_inst.traffic_state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _151_ (.CLK(net13),
    .D(_017_),
    .RESET_B(net11),
    .Q(\mod.traffic_sm_inst.traffic_state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _152_ (.CLK(net12),
    .D(_001_),
    .RESET_B(net10),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[0] ));
 sky130_fd_sc_hd__dfrtp_1 _153_ (.CLK(net13),
    .D(_002_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[1] ));
 sky130_fd_sc_hd__dfrtp_1 _154_ (.CLK(net13),
    .D(_003_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[2] ));
 sky130_fd_sc_hd__dfrtp_1 _155_ (.CLK(net13),
    .D(_004_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[3] ));
 sky130_fd_sc_hd__dfrtp_1 _156_ (.CLK(net12),
    .D(_005_),
    .RESET_B(net10),
    .Q(\mod.cnter_enb_ovf_i1.cnt_val[4] ));
 sky130_fd_sc_hd__dfrtp_2 _157_ (.CLK(net13),
    .D(_000_),
    .RESET_B(net11),
    .Q(\mod.cnter_enb_ovf_i1.overflow ));
 sky130_fd_sc_hd__conb_1 tiny_user_project_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 tiny_user_project_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 tiny_user_project_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 tiny_user_project_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 tiny_user_project_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 tiny_user_project_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 tiny_user_project_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 tiny_user_project_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 tiny_user_project_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 tiny_user_project_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 tiny_user_project_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 tiny_user_project_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 tiny_user_project_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 tiny_user_project_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 tiny_user_project_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 tiny_user_project_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 tiny_user_project_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 tiny_user_project_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 tiny_user_project_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 tiny_user_project_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 tiny_user_project_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 tiny_user_project_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 tiny_user_project_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 tiny_user_project_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 tiny_user_project_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 tiny_user_project_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 tiny_user_project_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 tiny_user_project_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 tiny_user_project_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 tiny_user_project_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 tiny_user_project_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 tiny_user_project_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 tiny_user_project_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 tiny_user_project_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 tiny_user_project_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 tiny_user_project_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 tiny_user_project_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 tiny_user_project_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 tiny_user_project_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 tiny_user_project_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 tiny_user_project_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 tiny_user_project_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 tiny_user_project_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 tiny_user_project_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tiny_user_project_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tiny_user_project_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tiny_user_project_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tiny_user_project_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tiny_user_project_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tiny_user_project_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tiny_user_project_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tiny_user_project_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tiny_user_project_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tiny_user_project_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tiny_user_project_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 tiny_user_project_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 tiny_user_project_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 tiny_user_project_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 tiny_user_project_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 tiny_user_project_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 tiny_user_project_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 tiny_user_project_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 tiny_user_project_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 tiny_user_project_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 tiny_user_project_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 tiny_user_project_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 tiny_user_project_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 tiny_user_project_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 tiny_user_project_83 (.LO(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[10]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[10]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[8]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[9]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(io_out[21]));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(net3),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net2),
    .X(net13));
 sky130_fd_sc_hd__conb_1 tiny_user_project_14 (.LO(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(net2));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_188 ();
 assign io_oeb[0] = net14;
 assign io_oeb[10] = net24;
 assign io_oeb[11] = net25;
 assign io_oeb[12] = net26;
 assign io_oeb[13] = net27;
 assign io_oeb[14] = net28;
 assign io_oeb[15] = net29;
 assign io_oeb[16] = net30;
 assign io_oeb[17] = net31;
 assign io_oeb[18] = net32;
 assign io_oeb[19] = net33;
 assign io_oeb[1] = net15;
 assign io_oeb[20] = net34;
 assign io_oeb[21] = net35;
 assign io_oeb[22] = net36;
 assign io_oeb[23] = net37;
 assign io_oeb[24] = net38;
 assign io_oeb[25] = net39;
 assign io_oeb[26] = net40;
 assign io_oeb[27] = net41;
 assign io_oeb[28] = net42;
 assign io_oeb[29] = net43;
 assign io_oeb[2] = net16;
 assign io_oeb[30] = net44;
 assign io_oeb[31] = net45;
 assign io_oeb[32] = net46;
 assign io_oeb[33] = net47;
 assign io_oeb[34] = net48;
 assign io_oeb[35] = net49;
 assign io_oeb[36] = net50;
 assign io_oeb[37] = net51;
 assign io_oeb[3] = net17;
 assign io_oeb[4] = net18;
 assign io_oeb[5] = net19;
 assign io_oeb[6] = net20;
 assign io_oeb[7] = net21;
 assign io_oeb[8] = net22;
 assign io_oeb[9] = net23;
 assign io_out[0] = net52;
 assign io_out[10] = net62;
 assign io_out[11] = net63;
 assign io_out[12] = net64;
 assign io_out[13] = net65;
 assign io_out[14] = net66;
 assign io_out[15] = net67;
 assign io_out[1] = net53;
 assign io_out[22] = net68;
 assign io_out[23] = net69;
 assign io_out[24] = net70;
 assign io_out[25] = net71;
 assign io_out[26] = net72;
 assign io_out[27] = net73;
 assign io_out[28] = net74;
 assign io_out[29] = net75;
 assign io_out[2] = net54;
 assign io_out[30] = net76;
 assign io_out[31] = net77;
 assign io_out[32] = net78;
 assign io_out[33] = net79;
 assign io_out[34] = net80;
 assign io_out[35] = net81;
 assign io_out[36] = net82;
 assign io_out[37] = net83;
 assign io_out[3] = net55;
 assign io_out[4] = net56;
 assign io_out[5] = net57;
 assign io_out[6] = net58;
 assign io_out[7] = net59;
 assign io_out[8] = net60;
 assign io_out[9] = net61;
endmodule

