magic
tech sky130A
magscale 1 2
timestamp 1671710124
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 382 2128 19306 17876
<< metal2 >>
rect 386 19200 442 20000
rect 1122 19200 1178 20000
rect 1858 19200 1914 20000
rect 2594 19200 2650 20000
rect 3330 19200 3386 20000
rect 4066 19200 4122 20000
rect 4802 19200 4858 20000
rect 5538 19200 5594 20000
rect 6274 19200 6330 20000
rect 7010 19200 7066 20000
rect 7746 19200 7802 20000
rect 8482 19200 8538 20000
rect 9218 19200 9274 20000
rect 9954 19200 10010 20000
rect 10690 19200 10746 20000
rect 11426 19200 11482 20000
rect 12162 19200 12218 20000
rect 12898 19200 12954 20000
rect 13634 19200 13690 20000
rect 14370 19200 14426 20000
rect 15106 19200 15162 20000
rect 15842 19200 15898 20000
rect 16578 19200 16634 20000
rect 17314 19200 17370 20000
rect 18050 19200 18106 20000
rect 18786 19200 18842 20000
rect 19522 19200 19578 20000
<< obsm2 >>
rect 498 19144 1066 19258
rect 1234 19144 1802 19258
rect 1970 19144 2538 19258
rect 2706 19144 3274 19258
rect 3442 19144 4010 19258
rect 4178 19144 4746 19258
rect 4914 19144 5482 19258
rect 5650 19144 6218 19258
rect 6386 19144 6954 19258
rect 7122 19144 7690 19258
rect 7858 19144 8426 19258
rect 8594 19144 9162 19258
rect 9330 19144 9898 19258
rect 10066 19144 10634 19258
rect 10802 19144 11370 19258
rect 11538 19144 12106 19258
rect 12274 19144 12842 19258
rect 13010 19144 13578 19258
rect 13746 19144 14314 19258
rect 14482 19144 15050 19258
rect 15218 19144 15786 19258
rect 15954 19144 16522 19258
rect 16690 19144 17258 19258
rect 17426 19144 17994 19258
rect 18162 19144 18730 19258
rect 18898 19144 19300 19258
rect 388 1391 19300 19144
<< metal3 >>
rect 19200 18912 20000 19032
rect 19200 18504 20000 18624
rect 0 18232 800 18352
rect 19200 18096 20000 18216
rect 0 17824 800 17944
rect 19200 17688 20000 17808
rect 0 17416 800 17536
rect 19200 17280 20000 17400
rect 0 17008 800 17128
rect 19200 16872 20000 16992
rect 0 16600 800 16720
rect 19200 16464 20000 16584
rect 0 16192 800 16312
rect 19200 16056 20000 16176
rect 0 15784 800 15904
rect 19200 15648 20000 15768
rect 0 15376 800 15496
rect 19200 15240 20000 15360
rect 0 14968 800 15088
rect 19200 14832 20000 14952
rect 0 14560 800 14680
rect 19200 14424 20000 14544
rect 0 14152 800 14272
rect 19200 14016 20000 14136
rect 0 13744 800 13864
rect 19200 13608 20000 13728
rect 0 13336 800 13456
rect 19200 13200 20000 13320
rect 0 12928 800 13048
rect 19200 12792 20000 12912
rect 0 12520 800 12640
rect 19200 12384 20000 12504
rect 0 12112 800 12232
rect 19200 11976 20000 12096
rect 0 11704 800 11824
rect 19200 11568 20000 11688
rect 0 11296 800 11416
rect 19200 11160 20000 11280
rect 0 10888 800 11008
rect 19200 10752 20000 10872
rect 0 10480 800 10600
rect 19200 10344 20000 10464
rect 0 10072 800 10192
rect 19200 9936 20000 10056
rect 0 9664 800 9784
rect 19200 9528 20000 9648
rect 0 9256 800 9376
rect 19200 9120 20000 9240
rect 0 8848 800 8968
rect 19200 8712 20000 8832
rect 0 8440 800 8560
rect 19200 8304 20000 8424
rect 0 8032 800 8152
rect 19200 7896 20000 8016
rect 0 7624 800 7744
rect 19200 7488 20000 7608
rect 0 7216 800 7336
rect 19200 7080 20000 7200
rect 0 6808 800 6928
rect 19200 6672 20000 6792
rect 0 6400 800 6520
rect 19200 6264 20000 6384
rect 0 5992 800 6112
rect 19200 5856 20000 5976
rect 0 5584 800 5704
rect 19200 5448 20000 5568
rect 0 5176 800 5296
rect 19200 5040 20000 5160
rect 0 4768 800 4888
rect 19200 4632 20000 4752
rect 0 4360 800 4480
rect 19200 4224 20000 4344
rect 0 3952 800 4072
rect 19200 3816 20000 3936
rect 0 3544 800 3664
rect 19200 3408 20000 3528
rect 0 3136 800 3256
rect 19200 3000 20000 3120
rect 0 2728 800 2848
rect 19200 2592 20000 2712
rect 0 2320 800 2440
rect 19200 2184 20000 2304
rect 0 1912 800 2032
rect 19200 1776 20000 1896
rect 0 1504 800 1624
rect 19200 1368 20000 1488
rect 19200 960 20000 1080
<< obsm3 >>
rect 800 18832 19120 19005
rect 800 18704 19212 18832
rect 800 18432 19120 18704
rect 880 18424 19120 18432
rect 880 18296 19212 18424
rect 880 18152 19120 18296
rect 800 18024 19120 18152
rect 880 18016 19120 18024
rect 880 17888 19212 18016
rect 880 17744 19120 17888
rect 800 17616 19120 17744
rect 880 17608 19120 17616
rect 880 17480 19212 17608
rect 880 17336 19120 17480
rect 800 17208 19120 17336
rect 880 17200 19120 17208
rect 880 17072 19212 17200
rect 880 16928 19120 17072
rect 800 16800 19120 16928
rect 880 16792 19120 16800
rect 880 16664 19212 16792
rect 880 16520 19120 16664
rect 800 16392 19120 16520
rect 880 16384 19120 16392
rect 880 16256 19212 16384
rect 880 16112 19120 16256
rect 800 15984 19120 16112
rect 880 15976 19120 15984
rect 880 15848 19212 15976
rect 880 15704 19120 15848
rect 800 15576 19120 15704
rect 880 15568 19120 15576
rect 880 15440 19212 15568
rect 880 15296 19120 15440
rect 800 15168 19120 15296
rect 880 15160 19120 15168
rect 880 15032 19212 15160
rect 880 14888 19120 15032
rect 800 14760 19120 14888
rect 880 14752 19120 14760
rect 880 14624 19212 14752
rect 880 14480 19120 14624
rect 800 14352 19120 14480
rect 880 14344 19120 14352
rect 880 14216 19212 14344
rect 880 14072 19120 14216
rect 800 13944 19120 14072
rect 880 13936 19120 13944
rect 880 13808 19212 13936
rect 880 13664 19120 13808
rect 800 13536 19120 13664
rect 880 13528 19120 13536
rect 880 13400 19212 13528
rect 880 13256 19120 13400
rect 800 13128 19120 13256
rect 880 13120 19120 13128
rect 880 12992 19212 13120
rect 880 12848 19120 12992
rect 800 12720 19120 12848
rect 880 12712 19120 12720
rect 880 12584 19212 12712
rect 880 12440 19120 12584
rect 800 12312 19120 12440
rect 880 12304 19120 12312
rect 880 12176 19212 12304
rect 880 12032 19120 12176
rect 800 11904 19120 12032
rect 880 11896 19120 11904
rect 880 11768 19212 11896
rect 880 11624 19120 11768
rect 800 11496 19120 11624
rect 880 11488 19120 11496
rect 880 11360 19212 11488
rect 880 11216 19120 11360
rect 800 11088 19120 11216
rect 880 11080 19120 11088
rect 880 10952 19212 11080
rect 880 10808 19120 10952
rect 800 10680 19120 10808
rect 880 10672 19120 10680
rect 880 10544 19212 10672
rect 880 10400 19120 10544
rect 800 10272 19120 10400
rect 880 10264 19120 10272
rect 880 10136 19212 10264
rect 880 9992 19120 10136
rect 800 9864 19120 9992
rect 880 9856 19120 9864
rect 880 9728 19212 9856
rect 880 9584 19120 9728
rect 800 9456 19120 9584
rect 880 9448 19120 9456
rect 880 9320 19212 9448
rect 880 9176 19120 9320
rect 800 9048 19120 9176
rect 880 9040 19120 9048
rect 880 8912 19212 9040
rect 880 8768 19120 8912
rect 800 8640 19120 8768
rect 880 8632 19120 8640
rect 880 8504 19212 8632
rect 880 8360 19120 8504
rect 800 8232 19120 8360
rect 880 8224 19120 8232
rect 880 8096 19212 8224
rect 880 7952 19120 8096
rect 800 7824 19120 7952
rect 880 7816 19120 7824
rect 880 7688 19212 7816
rect 880 7544 19120 7688
rect 800 7416 19120 7544
rect 880 7408 19120 7416
rect 880 7280 19212 7408
rect 880 7136 19120 7280
rect 800 7008 19120 7136
rect 880 7000 19120 7008
rect 880 6872 19212 7000
rect 880 6728 19120 6872
rect 800 6600 19120 6728
rect 880 6592 19120 6600
rect 880 6464 19212 6592
rect 880 6320 19120 6464
rect 800 6192 19120 6320
rect 880 6184 19120 6192
rect 880 6056 19212 6184
rect 880 5912 19120 6056
rect 800 5784 19120 5912
rect 880 5776 19120 5784
rect 880 5648 19212 5776
rect 880 5504 19120 5648
rect 800 5376 19120 5504
rect 880 5368 19120 5376
rect 880 5240 19212 5368
rect 880 5096 19120 5240
rect 800 4968 19120 5096
rect 880 4960 19120 4968
rect 880 4832 19212 4960
rect 880 4688 19120 4832
rect 800 4560 19120 4688
rect 880 4552 19120 4560
rect 880 4424 19212 4552
rect 880 4280 19120 4424
rect 800 4152 19120 4280
rect 880 4144 19120 4152
rect 880 4016 19212 4144
rect 880 3872 19120 4016
rect 800 3744 19120 3872
rect 880 3736 19120 3744
rect 880 3608 19212 3736
rect 880 3464 19120 3608
rect 800 3336 19120 3464
rect 880 3328 19120 3336
rect 880 3200 19212 3328
rect 880 3056 19120 3200
rect 800 2928 19120 3056
rect 880 2920 19120 2928
rect 880 2792 19212 2920
rect 880 2648 19120 2792
rect 800 2520 19120 2648
rect 880 2512 19120 2520
rect 880 2384 19212 2512
rect 880 2240 19120 2384
rect 800 2112 19120 2240
rect 880 2104 19120 2112
rect 880 1976 19212 2104
rect 880 1832 19120 1976
rect 800 1704 19120 1832
rect 880 1696 19120 1704
rect 880 1568 19212 1696
rect 880 1424 19120 1568
rect 800 1395 19120 1424
<< metal4 >>
rect 3163 2128 3483 17456
rect 5382 2128 5702 17456
rect 7602 2128 7922 17456
rect 9821 2128 10141 17456
rect 12041 2128 12361 17456
rect 14260 2128 14580 17456
rect 16480 2128 16800 17456
rect 18699 2128 19019 17456
<< obsm4 >>
rect 10547 17536 17053 18597
rect 10547 8467 11961 17536
rect 12441 8467 14180 17536
rect 14660 8467 16400 17536
rect 16880 8467 17053 17536
<< labels >>
rlabel metal3 s 19200 960 20000 1080 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 19200 13200 20000 13320 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 19200 14424 20000 14544 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 19200 15648 20000 15768 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 19200 16872 20000 16992 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 19200 18096 20000 18216 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 19522 19200 19578 20000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 17314 19200 17370 20000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 15106 19200 15162 20000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 12898 19200 12954 20000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 10690 19200 10746 20000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 8482 19200 8538 20000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 6274 19200 6330 20000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 4066 19200 4122 20000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 1858 19200 1914 20000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 19200 3408 20000 3528 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 19200 4632 20000 4752 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 19200 5856 20000 5976 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 19200 7080 20000 7200 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 19200 8304 20000 8424 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 19200 11976 20000 12096 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 19200 1776 20000 1896 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 19200 14016 20000 14136 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 19200 15240 20000 15360 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 19200 16464 20000 16584 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 19200 17688 20000 17808 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 19200 18912 20000 19032 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 18050 19200 18106 20000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 15842 19200 15898 20000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 13634 19200 13690 20000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 11426 19200 11482 20000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 9218 19200 9274 20000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 19200 3000 20000 3120 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 7010 19200 7066 20000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 4802 19200 4858 20000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 2594 19200 2650 20000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 386 19200 442 20000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 19200 4224 20000 4344 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 19200 5448 20000 5568 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 19200 6672 20000 6792 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 19200 7896 20000 8016 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 19200 9120 20000 9240 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 19200 10344 20000 10464 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 19200 11568 20000 11688 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 19200 12792 20000 12912 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 19200 1368 20000 1488 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 19200 13608 20000 13728 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 19200 14832 20000 14952 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 19200 16056 20000 16176 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 19200 17280 20000 17400 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 19200 18504 20000 18624 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 18786 19200 18842 20000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 16578 19200 16634 20000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 14370 19200 14426 20000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 12162 19200 12218 20000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 9954 19200 10010 20000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 19200 2592 20000 2712 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 7746 19200 7802 20000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 5538 19200 5594 20000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 3330 19200 3386 20000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 1122 19200 1178 20000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 19200 3816 20000 3936 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 1912 800 2032 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 19200 5040 20000 5160 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 19200 6264 20000 6384 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 19200 7488 20000 7608 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 19200 8712 20000 8832 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 19200 9936 20000 10056 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 19200 11160 20000 11280 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 19200 12384 20000 12504 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 3163 2128 3483 17456 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 17456 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 17456 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 17456 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 5382 2128 5702 17456 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 9821 2128 10141 17456 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 14260 2128 14580 17456 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 18699 2128 19019 17456 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 875908
string GDS_FILE /home/runner/work/traffic_controller/traffic_controller/openlane/tiny_user_project/runs/22_12_22_11_53/results/signoff/tiny_user_project.magic.gds
string GDS_START 286188
<< end >>

